@00000000
97 21 00 00 93 81 41 87 17 01 02 00 13 01 81 FF
33 04 01 00 6F 00 40 00
@00000018
13 01 01 FE 23 2E 81 00 13 04 01 02 93 07 40 00
23 26 F4 FE 93 07 C0 00 23 24 F4 FE 03 27 C4 FE
83 27 84 FE B3 07 F7 00 23 22 F4 FE 6F F0 1F FF
@00000048
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
98 FF FF FF 18 00 00 00 00 00 00 00
