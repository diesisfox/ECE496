@00000000
97 11 00 00 93 81 C1 07 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 C0 7A
@00000018
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 83 25 C4 FE 13 88 05 00 93 D5 F5 41
93 88 05 00 83 25 84 FE 13 86 05 00 93 D5 F5 41
93 86 05 00 33 85 C8 02 B3 85 06 03 B3 05 B5 00
33 05 C8 02 B3 37 C8 02 13 07 05 00 B3 86 F5 00
93 87 06 00 93 96 67 00 13 53 A7 01 33 E3 66 00
93 D3 A7 41 93 07 03 00 13 85 07 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 03 C7 C1 80 93 07 20 01 63 08 F7 08
83 C7 C1 80 93 86 07 00 B7 17 00 00 13 87 47 80
93 97 26 00 B3 07 F7 00 83 A7 07 00 23 26 F4 FE
03 27 C4 FE 93 07 07 00 93 97 27 00 B3 87 E7 00
93 97 57 00 13 87 07 00 B7 17 00 00 83 A7 C7 87
33 07 F7 00 B7 17 00 00 23 AE E7 86 03 27 C4 FE
93 07 07 00 93 97 47 00 B3 87 E7 40 93 97 37 00
13 87 07 00 B7 17 00 00 83 A7 07 88 33 07 F7 00
B7 17 00 00 23 A0 E7 88 83 C7 C1 80 93 87 17 00
13 F7 F7 0F 23 86 E1 80 6F 00 80 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 83 C7 C1 80 63 82 07 1A
83 C7 C1 80 93 87 F7 FF 13 F7 F7 0F 23 86 E1 80
83 C7 C1 80 63 94 07 02 B7 17 00 00 37 A7 03 FA
13 07 A7 99 23 AE E7 86 B7 17 00 00 37 A7 A3 FC
13 07 A7 99 23 A0 E7 88 6F 00 C0 16 83 C7 C1 80
93 86 07 00 B7 17 00 00 13 87 47 80 93 97 26 00
B3 07 F7 00 83 A7 07 00 23 26 F4 FE 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 57 00
33 07 F0 40 B7 17 00 00 83 A7 C7 87 33 07 F7 00
B7 17 00 00 23 AE E7 86 03 27 C4 FE 93 07 07 00
13 17 47 00 B3 87 E7 40 93 97 37 00 13 87 07 00
B7 17 00 00 83 A7 07 88 33 07 F7 00 B7 17 00 00
23 A0 E7 88 03 27 C4 FE 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 77 00 33 87 E7 40 B7 17 00 00
83 A7 C7 87 33 07 F7 00 B7 67 FC 02 93 87 67 66
63 D2 E7 02 03 27 C4 FE 93 07 10 D8 33 07 F7 02
B7 67 FC 02 93 87 67 66 33 07 F7 00 B7 17 00 00
23 AE E7 86 03 27 C4 FE 93 07 07 00 93 97 47 00
B3 87 E7 40 93 97 57 00 33 87 E7 40 B7 17 00 00
83 A7 07 88 33 07 F7 00 B7 67 5C 03 93 87 67 66
63 D2 E7 02 03 27 C4 FE 93 07 10 E2 33 07 F7 02
B7 67 5C 03 93 87 67 66 33 07 F7 00 B7 17 00 00
23 A0 E7 88 B7 17 00 00 03 A7 C7 87 B7 A7 03 FA
93 87 A7 99 63 5A F7 00 B7 17 00 00 37 A7 03 FA
13 07 A7 99 23 AE E7 86 B7 17 00 00 03 A7 07 88
B7 A7 A3 FC 93 87 A7 99 63 5E F7 00 B7 17 00 00
37 A7 A3 FC 13 07 A7 99 23 A0 E7 88 6F 00 80 00
13 00 00 00 03 24 C1 01 13 01 01 02 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
A3 0F F4 FC 83 C7 C1 80 93 86 07 00 B7 17 00 00
13 87 47 80 93 97 26 00 B3 07 F7 00 83 A7 07 00
23 26 F4 FE 83 47 F4 FD 93 F7 27 00 63 82 07 02
83 27 C4 FE 13 97 67 00 B7 17 00 00 83 A7 07 88
33 07 F7 00 B7 17 00 00 23 A0 E7 88 6F 00 C0 02
83 47 F4 FD 93 F7 47 00 63 80 07 02 B7 17 00 00
03 A7 07 88 83 27 C4 FE 93 97 67 00 33 07 F7 40
B7 17 00 00 23 A0 E7 88 83 47 F4 FD 93 F7 17 00
63 82 07 02 83 27 C4 FE 13 97 67 00 B7 17 00 00
83 A7 C7 87 33 07 F7 00 B7 17 00 00 23 AE E7 86
6F 00 C0 02 83 47 F4 FD 93 F7 87 00 63 80 07 02
B7 17 00 00 03 A7 C7 87 83 27 C4 FE 93 97 67 00
33 07 F7 40 B7 17 00 00 23 AE E7 86 03 27 C4 FE
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 77 00
33 87 E7 40 B7 17 00 00 83 A7 C7 87 33 07 F7 00
B7 67 FC 02 93 87 67 66 63 D2 E7 02 03 27 C4 FE
93 07 10 D8 33 07 F7 02 B7 67 FC 02 93 87 67 66
33 07 F7 00 B7 17 00 00 23 AE E7 86 03 27 C4 FE
93 07 07 00 93 97 47 00 B3 87 E7 40 93 97 57 00
33 87 E7 40 B7 17 00 00 83 A7 07 88 33 07 F7 00
B7 67 5C 03 93 87 67 66 63 D2 E7 02 03 27 C4 FE
93 07 10 E2 33 07 F7 02 B7 67 5C 03 93 87 67 66
33 07 F7 00 B7 17 00 00 23 A0 E7 88 B7 17 00 00
03 A7 C7 87 B7 A7 03 FA 93 87 A7 99 63 5A F7 00
B7 17 00 00 37 A7 03 FA 13 07 A7 99 23 AE E7 86
B7 17 00 00 03 A7 07 88 B7 A7 A3 FC 93 87 A7 99
63 5A F7 00 B7 17 00 00 37 A7 A3 FC 13 07 A7 99
23 A0 E7 88 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FC 23 2E 11 02 23 2C 81 02
13 04 01 04 23 26 A4 FC 23 24 B4 FC 93 07 F0 0F
23 12 F4 FE 23 26 04 FE 23 24 04 FE 23 13 04 FE
6F 00 C0 08 83 25 C4 FE 03 25 C4 FE EF F0 5F B0
23 20 A4 FE 83 25 84 FE 03 25 84 FE EF F0 5F AF
23 2E A4 FC 03 27 04 FE 83 27 C4 FD 33 07 F7 00
B7 07 00 10 63 C4 E7 06 03 27 04 FE 83 27 C4 FD
B3 07 F7 40 03 27 C4 FC B3 07 F7 00 23 2C F4 FC
83 25 84 FE 03 25 C4 FE EF F0 9F AB 93 07 05 00
93 97 17 00 03 27 84 FC B3 07 F7 00 23 2A F4 FC
83 27 84 FD 23 26 F4 FE 83 27 44 FD 23 24 F4 FE
83 57 64 FE 93 87 17 00 23 13 F4 FE 03 57 64 FE
83 57 44 FE E3 F8 E7 F6 6F 00 80 00 13 00 00 00
83 57 64 FE 93 F7 F7 0F 13 85 07 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 83 C7 C1 80
93 86 07 00 B7 17 00 00 13 87 47 80 93 97 26 00
B3 07 F7 00 83 A7 07 00 23 2E F4 FC B7 17 00 00
83 A7 07 88 23 26 F4 FE 23 24 04 FE 6F 00 00 08
B7 17 00 00 83 A7 C7 87 23 22 F4 FE 23 20 04 FE
6F 00 40 04 83 25 C4 FE 03 25 44 FE EF F0 9F EB
93 07 05 00 A3 0D F4 FC B7 17 00 00 83 A7 47 88
03 47 B4 FD 23 A6 E7 00 03 27 44 FE 83 27 C4 FD
B3 07 F7 00 23 22 F4 FE 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 93 07 F0 27 E3 FC E7 FA
03 27 C4 FE 83 27 C4 FD B3 07 F7 00 23 26 F4 FE
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
93 07 F0 1D E3 FE E7 F6 13 00 00 00 13 00 00 00
83 20 C1 02 03 24 81 02 13 01 01 03 67 80 00 00
13 01 01 FE 23 2E 81 00 13 04 01 02 B7 17 00 00
83 A7 47 88 23 A8 07 00 23 26 04 FE 6F 00 00 05
13 07 F0 0F 83 27 C4 FE B3 07 F7 40 13 97 07 01
93 06 F0 0F 83 27 C4 FE B3 87 F6 40 93 97 87 00
B3 66 F7 00 13 07 F0 0F 83 27 C4 FE 33 07 F7 40
B7 17 00 00 83 A7 47 88 33 E7 E6 00 23 AA E7 00
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
93 07 E0 0F E3 F6 E7 FA 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 B7 17 00 00 83 A7 47 88
23 A8 07 00 23 26 04 FE 6F 00 00 05 13 07 F0 0F
83 27 C4 FE B3 07 F7 40 13 97 07 01 93 06 F0 0F
83 27 C4 FE B3 87 F6 40 93 97 87 00 B3 66 F7 00
13 07 F0 0F 83 27 C4 FE 33 07 F7 40 B7 17 00 00
83 A7 47 88 33 E7 E6 00 23 AA E7 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 E0 0F
E3 F6 E7 FA 13 00 00 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FF 23 26 11 00
23 24 81 00 13 04 01 01 B7 17 00 00 83 A7 47 88
13 07 10 00 23 A0 E7 00 EF F0 9F EC B7 17 00 00
83 A7 47 88 23 A2 07 00 B7 17 00 00 83 A7 47 88
23 A4 07 00 EF F0 9F DC 6F 00 00 00
@00000804
9A 99 03 00 CD CC 01 00 66 E6 00 00 33 73 00 00
9A 39 00 00 CD 1C 00 00 66 0E 00 00 33 07 00 00
9A 03 00 00 CD 01 00 00 E6 00 00 00 73 00 00 00
3A 00 00 00 1D 00 00 00 0E 00 00 00 07 00 00 00
04 00 00 00 02 00 00 00 01 00 00 00
@00000850
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
90 F7 FF FF 18 00 00 00 00 00 00 00
@0000087C
9A 99 03 FA 9A 99 A3 FC 00 00 00 80
