@00000000
97 31 00 00 93 81 81 48 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 40 00
@00000018
B7 37 00 00 03 A6 C7 C8 13 01 01 FF B7 17 00 00
93 87 07 BF 23 26 11 00 13 07 10 00 93 85 C7 06
23 20 E6 00 93 87 87 46 83 A6 07 00 13 87 07 00
93 87 C7 FF 23 2A D6 00 E3 98 E5 FE EF 00 C0 6B
E3 1E 05 FE EF 00 C0 50 E3 1A 05 FE EF 00 40 50
E3 0A 05 FE 6F F0 9F FE B3 07 B5 02 33 15 B5 02
93 D7 A7 01 13 15 65 00 33 65 F5 00 67 80 00 00
83 C6 41 81 93 07 20 01 63 8A F6 04 B7 17 00 00
13 97 26 00 93 87 07 BF B3 87 E7 00 03 A6 07 00
37 35 00 00 03 A3 C1 80 83 28 05 C9 13 17 26 00
93 17 46 00 33 07 C7 00 B3 87 C7 40 13 17 57 00
93 97 37 00 33 07 67 00 B3 87 17 01 93 86 16 00
23 A6 E1 80 23 28 F5 C8 23 8A D1 80 67 80 00 00
83 C7 41 81 63 88 07 0C 93 87 F7 FF 93 F7 F7 0F
23 8A F1 80 63 82 07 0C 37 17 00 00 13 07 07 BF
93 97 27 00 B3 07 F7 00 83 A6 07 00 37 38 00 00
03 25 08 C9 83 A5 C1 80 13 97 26 00 93 97 46 00
33 07 D7 00 33 86 F6 40 13 13 57 00 13 16 36 00
13 17 77 00 B3 85 65 40 33 06 A6 00 33 07 D7 40
37 65 FC 02 23 A6 B1 80 23 28 C8 C8 33 07 B7 00
13 05 65 66 63 5A E5 00 93 05 10 D8 B3 85 B6 02
B3 85 A5 00 23 A6 B1 80 B3 87 D7 40 93 97 57 00
B3 87 D7 40 37 67 5C 03 B3 87 C7 00 13 07 67 66
63 5A F7 00 93 07 10 E2 B3 86 F6 02 33 86 E6 00
23 28 C8 C8 B7 A7 03 FA 93 87 A7 99 63 D4 F5 00
23 A6 F1 80 B7 A7 A3 FC 93 87 A7 99 63 54 F6 00
23 28 F8 C8 67 80 00 00 B7 A7 03 FA 93 87 A7 99
23 A6 F1 80 B7 A7 A3 FC 37 37 00 00 93 87 A7 99
23 28 F7 C8 67 80 00 00 83 C7 41 81 B7 35 00 00
03 A8 05 C9 13 97 27 00 B7 17 00 00 93 87 07 BF
B3 87 E7 00 13 77 25 00 83 A7 07 00 63 02 07 0C
13 97 67 00 33 08 E8 00 23 A8 05 C9 13 77 15 00
83 A6 C1 80 63 0A 07 08 13 97 67 00 B3 86 E6 00
23 A6 D1 80 13 97 27 00 33 07 F7 00 13 17 77 00
33 07 F7 40 37 66 FC 02 33 07 D7 00 13 06 66 66
63 5A E6 00 93 06 10 D8 B3 86 D7 02 B3 86 C6 00
23 A6 D1 80 13 97 47 00 33 07 F7 40 13 17 57 00
33 07 F7 40 37 66 5C 03 33 07 07 01 13 06 66 66
63 5A E6 00 13 07 10 E2 B3 87 E7 02 33 88 C7 00
23 A8 05 C9 37 A7 03 FA 13 07 A7 99 63 D4 E6 00
23 A6 E1 80 37 A7 A3 FC 13 07 A7 99 63 54 E8 00
23 A8 E5 C8 67 80 00 00 13 75 85 00 E3 0C 05 F6
13 97 67 00 B3 86 E6 40 23 A6 D1 80 6F F0 9F F6
13 77 45 00 E3 04 07 F4 13 97 67 00 33 08 E8 40
23 A8 05 C9 6F F0 9F F3 13 0E 05 00 13 03 00 00
13 07 00 00 13 06 00 00 93 0F 00 00 13 08 00 00
93 07 00 00 93 06 00 00 93 0E F0 0F 37 0F 00 10
B3 8F FF 02 13 03 13 00 33 07 07 41 13 13 03 01
33 07 C7 01 13 53 03 01 B3 86 C6 02 33 B5 C7 02
B3 86 F6 01 93 5F F7 41 B3 87 C7 02 B3 86 A6 00
93 96 66 00 13 06 07 00 93 D7 A7 01 B3 E7 F6 00
93 97 17 00 B3 87 B7 00 63 00 D3 05 33 05 C6 02
93 D6 F7 41 33 17 C6 02 13 55 A5 01 B3 88 F7 02
13 17 67 00 33 67 A7 00 33 98 F7 02 93 D8 A8 01
13 18 68 00 33 68 18 01 33 05 E8 00 E3 52 AF F8
13 75 F3 0F 67 80 00 00 13 05 F0 0F 67 80 00 00
83 C7 41 81 13 01 01 FF 23 26 81 00 13 97 27 00
B7 17 00 00 93 87 07 BF B3 87 E7 00 83 AF 07 00
B7 37 00 00 03 A3 07 C9 03 A4 C1 80 B7 37 00 00
83 A2 C7 C8 23 24 91 00 93 03 00 1E 13 0E F0 0F
B7 0E 00 10 93 08 04 00 13 0F 00 28 13 05 00 00
93 05 00 00 93 07 00 00 93 06 00 00 13 07 00 00
13 06 00 00 13 08 00 00 33 08 F8 02 33 07 B7 40
13 05 15 00 13 15 05 01 33 07 17 01 13 55 05 01
B3 86 C6 02 B3 B5 C7 02 B3 86 06 01 13 58 F7 41
B3 87 C7 02 B3 86 B6 00 93 96 66 00 13 06 07 00
93 D7 A7 01 B3 E7 F6 00 93 97 17 00 B3 87 67 00
63 02 C5 07 B3 05 C6 02 93 D6 F7 41 33 17 C6 02
93 D5 A5 01 13 17 67 00 33 67 B7 00 B3 84 F7 02
B3 95 F7 02 93 D4 A4 01 93 95 65 00 B3 E5 95 00
B3 04 B7 00 E3 D2 9E F8 23 A6 A2 00 13 0F FF FF
B3 88 F8 01 E3 1C 0F F4 93 83 F3 FF 33 03 F3 01
E3 92 03 F4 03 24 C1 00 83 24 81 00 13 01 01 01
67 80 00 00 13 05 F0 0F 23 A6 A2 00 13 0F FF FF
B3 88 F8 01 E3 14 0F F2 6F F0 1F FD 93 07 10 00
B3 96 D7 00 63 5E D0 02 B7 37 00 00 03 A7 C7 C8
13 08 00 00 B3 07 B8 00 23 24 F7 00 23 22 A7 00
93 07 00 00 93 87 17 00 23 26 C7 00 93 F7 F7 0F
E3 CA D7 FE 13 08 18 00 13 78 F8 0F E3 4C D8 FC
67 80 00 00 93 57 15 00 13 97 27 00 B7 17 00 00
93 87 07 BF B3 87 E7 00 13 75 15 00 37 37 00 00
83 A7 C7 04 83 26 C7 C8 63 0E 05 00 13 86 07 40
03 A7 07 00 93 87 47 00 23 AA E6 00 E3 1A F6 FE
67 80 00 00 13 87 C7 3F 83 25 07 00 13 06 07 00
13 07 C7 FF 23 AA B6 00 E3 98 C7 FE 67 80 00 00
B7 37 00 00 03 A7 87 C8 13 01 01 FF 23 20 21 01
23 22 91 00 83 A7 01 81 83 24 07 00 23 26 11 00
23 24 81 00 13 05 00 00 63 8C 97 08 93 C7 F7 FF
33 F4 97 00 93 77 F4 00 63 92 07 0A 93 77 04 01
63 82 07 06 83 C6 41 81 93 07 20 01 13 05 10 00
63 8A F6 04 B7 17 00 00 13 97 26 00 93 87 07 BF
B3 87 E7 00 03 A6 07 00 37 38 00 00 03 AE C1 80
03 23 08 C9 13 17 26 00 93 17 46 00 33 07 C7 00
B3 87 C7 40 13 17 57 00 93 97 37 00 33 07 C7 01
B3 87 67 00 93 86 16 00 23 A6 E1 80 23 28 F8 C8
23 8A D1 80 13 74 04 02 63 16 04 0A 83 A7 01 81
B3 C7 F4 00 93 D7 67 00 93 F7 F7 00 63 9C 07 02
83 20 C1 00 03 24 81 00 23 A8 91 80 83 24 41 00
03 29 01 00 13 01 01 01 67 80 00 00 13 85 07 00
EF F0 9F B9 93 77 04 01 13 05 10 00 E3 8C 07 FA
6F F0 5F F5 93 D7 64 00 93 F7 F7 0F 93 96 17 00
13 F7 C6 01 B7 16 00 00 93 86 06 BF B3 86 E6 00
13 F7 17 00 83 A7 C6 04 B7 36 00 00 83 A6 C6 C8
63 0A 07 04 13 86 07 40 03 A7 07 00 93 87 47 00
23 AA E6 00 E3 1A F6 FE 83 20 C1 00 03 24 81 00
23 A8 91 80 83 24 41 00 03 29 01 00 13 01 01 01
67 80 00 00 EF F0 DF A2 83 A7 01 81 13 05 10 00
B3 C7 F4 00 93 D7 67 00 93 F7 F7 00 E3 8A 07 F4
6F F0 5F F8 13 87 C7 3F 83 25 07 00 13 06 07 00
13 07 C7 FF 23 AA B6 00 E3 98 C7 FE 83 20 C1 00
03 24 81 00 23 A8 91 80 83 24 41 00 03 29 01 00
13 01 01 01 67 80 00 00 83 C7 41 81 13 01 01 FB
23 20 21 05 13 97 27 00 B7 17 00 00 93 87 07 BF
B3 87 E7 00 83 A7 07 00 37 37 00 00 03 29 07 C9
23 2C 41 03 23 28 61 03 23 26 71 03 23 24 81 03
23 26 11 04 23 24 81 04 23 22 91 04 23 2E 31 03
23 2A 51 03 23 22 91 03 23 20 A1 03 23 2E B1 01
23 20 F1 00 13 9C 57 00 13 0B 00 02 13 05 00 00
37 0A 00 10 B7 3B 00 00 83 A4 C1 80 13 0D 0B FE
93 0A 00 00 93 09 F0 0F B7 1C 00 00 13 04 00 00
13 06 00 00 93 07 00 00 13 08 00 00 13 07 00 00
93 06 00 00 93 05 00 00 B3 85 F5 02 33 07 C7 40
33 07 97 00 13 04 14 00 13 14 04 01 13 54 04 01
33 08 D8 02 33 B6 F6 02 B3 85 05 01 B3 87 F6 02
93 06 07 00 33 87 C5 00 13 17 67 00 93 D5 F6 41
93 D7 A7 01 B3 67 F7 00 93 97 17 00 B3 87 27 01
63 0E 34 37 33 86 D6 02 13 D8 F7 41 33 97 D6 02
13 56 A6 01 13 17 67 00 33 67 C7 00 B3 88 F7 02
33 96 F7 02 93 D8 A8 01 13 16 66 00 33 66 16 01
B3 08 C7 00 E3 52 1A F9 93 07 04 00 33 05 F5 00
63 C8 AC 2E 83 A7 CB C8 93 06 0D 00 23 A4 D7 00
23 A2 57 01 13 07 00 02 13 07 F7 FF 23 A6 87 00
13 77 F7 0F E3 1A 07 FE 93 86 16 00 E3 10 DB FE
93 8A 0A 02 13 07 00 28 B3 84 84 01 E3 90 EA F2
13 0B 0B 02 13 07 00 20 33 09 89 01 E3 1E EB EE
13 0C 40 00 93 09 F0 0F 37 0A 00 10 37 37 00 00
03 29 07 C9 03 27 01 00 93 05 00 00 93 08 00 1E
B3 1C 87 01 13 08 00 28 13 07 0C 00 13 04 10 00
B3 D8 88 41 33 58 88 41 33 14 84 01 13 9D 1C 00
13 8C 05 00 93 05 07 00 83 A4 C1 80 13 07 08 00
33 1B BC 00 93 7D 1C 00 13 08 0C 00 B3 84 9C 00
93 0A 10 00 37 13 00 00 13 0C 07 00 6F 00 C0 00
B3 04 9D 00 93 8A 1A 00 93 8E FA FF 33 E7 DD 01
B3 84 94 41 E3 06 07 FE 13 0E 00 00 93 06 00 00
13 07 00 00 93 0F 00 00 93 02 00 00 13 06 00 00
13 0F 00 00 33 0F EF 02 B3 86 D2 40 B3 86 96 00
13 0E 1E 00 13 1E 0E 01 13 5E 0E 01 B3 8F CF 02
B3 32 E6 02 33 0F FF 01 33 07 E6 02 13 86 06 00
B3 06 5F 00 93 96 66 00 13 5F F6 41 13 57 A7 01
33 E7 E6 00 13 17 17 00 33 07 27 01 63 0A 3E 23
B3 06 C6 02 93 5F F7 41 B3 12 C6 02 93 D6 A6 01
93 92 62 00 B3 E2 D2 00 B3 03 E7 02 B3 16 E7 02
93 D3 A3 01 93 96 66 00 B3 E6 76 00 B3 83 D2 00
E3 52 7A F8 93 06 0E 00 B3 9E BE 00 13 06 00 00
33 07 66 01 23 A4 E7 00 23 A2 D7 01 13 07 00 00
13 07 17 00 23 A6 D7 00 13 77 F7 0F E3 4A 87 FE
13 06 16 00 13 76 F6 0F E3 4C 86 FC 33 05 C5 01
63 4A A3 18 E3 E6 8A F1 13 07 0C 00 13 0C 08 00
13 0C 1C 00 13 08 07 00 33 09 99 01 E3 16 1C ED
13 8C F5 FF E3 14 0C E8 83 2C 01 00 37 37 00 00
83 24 07 C9 93 0A 00 00 13 0D 10 00 37 09 00 10
13 9B 1C 00 23 20 81 01 03 A4 C1 80 23 A4 57 01
93 FD 1A 00 33 04 94 01 13 0A 10 00 93 09 F0 0F
37 18 00 00 13 0C 00 28 6F 00 00 01 23 A2 A7 01
33 04 8B 00 13 0A 1A 00 13 07 FA FF 33 67 B7 01
33 04 94 41 E3 04 07 FE 93 06 00 00 93 0E 00 00
93 05 00 00 13 07 00 00 13 0E 00 00 13 06 00 00
13 03 00 00 33 03 E3 02 B3 86 DE 40 B3 86 86 00
93 85 15 00 93 95 05 01 93 D5 05 01 33 0E CE 02
B3 3E E6 02 33 03 C3 01 33 07 E6 02 13 86 06 00
B3 06 D3 01 93 96 66 00 13 53 F6 41 13 57 A7 01
33 E7 E6 00 13 17 17 00 33 07 97 00 63 84 35 11
B3 06 C6 02 13 5E F7 41 B3 1E C6 02 93 D6 A6 01
93 9E 6E 00 B3 EE DE 00 33 0F E7 02 B3 16 E7 02
13 5F AF 01 93 96 66 00 B3 E6 E6 01 33 8F DE 00
E3 52 E9 F9 13 87 05 00 33 05 B5 00 23 A6 E7 00
63 4E A8 08 63 04 8A 0B 83 A7 CB C8 6F F0 5F F3
EF F0 1F A4 E3 08 05 D0 13 0C 10 00 83 20 C1 04
03 24 81 04 83 24 41 04 03 29 01 04 83 29 C1 03
03 2A 81 03 83 2A 41 03 03 2B 01 03 83 2B C1 02
83 2C 41 02 03 2D 01 02 83 2D C1 01 13 05 0C 00
03 2C 81 02 13 01 01 05 67 80 00 00 93 07 F0 0F
6F F0 DF CB 23 26 B1 00 23 24 11 01 23 22 01 01
EF F0 1F 9E E3 12 05 FA 83 A7 CB C8 83 25 C1 00
83 28 81 00 03 28 41 00 37 13 00 00 6F F0 9F E4
93 06 F0 0F 13 0E F0 0F 6F F0 1F E0 EF F0 5F 9B
37 18 00 00 E3 1A 05 F6 E3 10 8A F7 93 8A 1A 00
93 07 00 1E B3 84 94 01 63 8C FA 00 83 A7 CB C8
6F F0 9F E5 13 07 F0 0F 93 05 F0 0F 6F F0 DF F2
03 2C 01 00 6F F0 9F F4
@00000BF0
9A 99 03 00 CD CC 01 00 66 E6 00 00 33 73 00 00
9A 39 00 00 CD 1C 00 00 66 0E 00 00 33 07 00 00
9A 03 00 00 CD 01 00 00 E6 00 00 00 73 00 00 00
3A 00 00 00 1D 00 00 00 0E 00 00 00 07 00 00 00
04 00 00 00 02 00 00 00 01 00 00 00 5C 10 00 00
5C 14 00 00 5C 18 00 00 5C 1C 00 00 5C 20 00 00
5C 24 00 00 5C 0C 00 00 5C 28 00 00 00 07 64 00
01 09 66 00 01 0A 67 00 02 0C 69 00 02 0D 6A 00
03 0F 6C 00 03 10 6E 00 04 12 6F 00 04 14 71 00
05 15 73 00 05 17 74 00 06 18 76 00 06 1A 77 00
07 1B 79 00 07 1D 7B 00 08 1F 7C 00 08 20 7E 00
09 22 7F 00 09 23 81 00 0A 25 83 00 0A 26 84 00
0B 28 86 00 0B 2A 88 00 0C 2B 89 00 0C 2D 8B 00
0D 2E 8C 00 0D 30 8E 00 0E 31 90 00 0E 33 91 00
0F 34 93 00 0F 36 94 00 10 38 96 00 10 39 98 00
11 3B 99 00 11 3C 9B 00 12 3E 9D 00 12 3F 9E 00
13 41 A0 00 13 43 A1 00 14 44 A3 00 14 46 A5 00
15 47 A6 00 15 49 A8 00 16 4A A9 00 16 4C AB 00
17 4E AD 00 17 4F AE 00 18 51 B0 00 18 52 B2 00
19 54 B3 00 19 55 B5 00 1A 57 B6 00 1A 59 B8 00
1B 5A BA 00 1B 5C BB 00 1C 5D BD 00 1C 5F BE 00
1D 60 C0 00 1D 62 C2 00 1E 64 C3 00 1E 65 C5 00
1F 67 C7 00 1F 68 C8 00 20 6A CA 00 21 6C CB 00
24 6E CC 00 27 70 CD 00 2A 73 CE 00 2E 75 CE 00
31 77 CF 00 34 7A D0 00 37 7C D1 00 3B 7E D2 00
3E 80 D3 00 41 83 D3 00 44 85 D4 00 47 87 D5 00
4B 8A D6 00 4E 8C D7 00 51 8E D7 00 54 91 D8 00
57 93 D9 00 5B 95 DA 00 5E 98 DB 00 61 9A DC 00
64 9C DC 00 68 9F DD 00 6B A1 DE 00 6E A3 DF 00
71 A6 E0 00 74 A8 E0 00 78 AA E1 00 7B AD E2 00
7E AF E3 00 81 B1 E4 00 84 B4 E4 00 88 B6 E5 00
8B B8 E6 00 8E BB E7 00 91 BD E8 00 95 BF E9 00
98 C1 E9 00 9B C4 EA 00 9E C6 EB 00 A1 C8 EC 00
A5 CB ED 00 A8 CD ED 00 AB CF EE 00 AE D2 EF 00
B2 D4 F0 00 B5 D6 F1 00 B8 D9 F2 00 BB DB F2 00
BE DD F3 00 C2 E0 F4 00 C5 E2 F5 00 C8 E4 F6 00
CB E7 F6 00 CE E9 F7 00 D2 EB F8 00 D5 EE F9 00
D8 F0 FA 00 DB F2 FB 00 DF F5 FB 00 E2 F7 FC 00
E5 F9 FD 00 E8 FC FE 00 EB FE FF 00 ED FE FD 00
ED FD F9 00 EE FC F5 00 EE FA F1 00 EE F9 ED 00
EF F8 E9 00 EF F6 E5 00 EF F5 E1 00 EF F4 DD 00
F0 F2 D9 00 F0 F1 D5 00 F0 F0 D1 00 F1 EE CD 00
F1 ED C9 00 F1 EC C5 00 F1 EA C1 00 F2 E9 BD 00
F2 E8 B9 00 F2 E6 B5 00 F3 E5 B1 00 F3 E4 AD 00
F3 E2 A9 00 F3 E1 A5 00 F4 E0 A1 00 F4 DE 9D 00
F4 DD 99 00 F4 DC 95 00 F5 DA 91 00 F5 D9 8D 00
F5 D8 89 00 F6 D6 85 00 F6 D5 81 00 F6 D4 7D 00
F6 D2 79 00 F7 D1 75 00 F7 D0 71 00 F7 CE 6D 00
F8 CD 69 00 F8 CC 65 00 F8 CA 61 00 F8 C9 5D 00
F9 C8 59 00 F9 C6 55 00 F9 C5 51 00 FA C4 4D 00
FA C2 49 00 FA C1 45 00 FA C0 41 00 FB BE 3D 00
FB BD 39 00 FB BC 35 00 FC BA 31 00 FC B9 2D 00
FC B8 29 00 FC B6 25 00 FD B5 21 00 FD B4 1D 00
FD B2 19 00 FE B1 15 00 FE B0 11 00 FE AE 0D 00
FE AD 09 00 FF AC 05 00 FF AA 01 00 FC A8 00 00
F8 A5 00 00 F4 A3 00 00 F0 A0 00 00 EC 9D 00 00
E8 9B 00 00 E4 98 00 00 E0 96 00 00 DC 93 00 00
D8 90 00 00 D4 8E 00 00 D0 8B 00 00 CC 88 00 00
C8 86 00 00 C4 83 00 00 C0 80 00 00 BC 7E 00 00
B8 7B 00 00 B4 79 00 00 B0 76 00 00 AC 73 00 00
A8 71 00 00 A4 6E 00 00 A0 6B 00 00 9C 69 00 00
98 66 00 00 94 64 00 00 90 61 00 00 8C 5E 00 00
88 5C 00 00 84 59 00 00 80 56 00 00 7C 54 00 00
78 51 00 00 74 4E 00 00 70 4C 00 00 6C 49 00 00
68 47 00 00 64 44 00 00 60 41 00 00 5C 3F 00 00
58 3C 00 00 54 39 00 00 50 37 00 00 4C 34 00 00
48 31 00 00 44 2F 00 00 40 2C 00 00 3C 2A 00 00
38 27 00 00 34 24 00 00 30 22 00 00 2C 1F 00 00
28 1C 00 00 24 1A 00 00 20 17 00 00 1C 14 00 00
18 12 00 00 14 0F 00 00 10 0D 00 00 0C 0A 00 00
08 07 00 00 04 05 00 00 00 02 00 00 FF FF FF 00
FE FE FE 00 FD FD FD 00 FC FC FC 00 FB FB FB 00
FA FA FA 00 F9 F9 F9 00 F8 F8 F8 00 F7 F7 F7 00
F6 F6 F6 00 F5 F5 F5 00 F4 F4 F4 00 F3 F3 F3 00
F2 F2 F2 00 F1 F1 F1 00 F0 F0 F0 00 EF EF EF 00
EE EE EE 00 ED ED ED 00 EC EC EC 00 EB EB EB 00
EA EA EA 00 E9 E9 E9 00 E8 E8 E8 00 E7 E7 E7 00
E6 E6 E6 00 E5 E5 E5 00 E4 E4 E4 00 E3 E3 E3 00
E2 E2 E2 00 E1 E1 E1 00 E0 E0 E0 00 DF DF DF 00
DE DE DE 00 DD DD DD 00 DC DC DC 00 DB DB DB 00
DA DA DA 00 D9 D9 D9 00 D8 D8 D8 00 D7 D7 D7 00
D6 D6 D6 00 D5 D5 D5 00 D4 D4 D4 00 D3 D3 D3 00
D2 D2 D2 00 D1 D1 D1 00 D0 D0 D0 00 CF CF CF 00
CE CE CE 00 CD CD CD 00 CC CC CC 00 CB CB CB 00
CA CA CA 00 C9 C9 C9 00 C8 C8 C8 00 C7 C7 C7 00
C6 C6 C6 00 C5 C5 C5 00 C4 C4 C4 00 C3 C3 C3 00
C2 C2 C2 00 C1 C1 C1 00 C0 C0 C0 00 BF BF BF 00
BE BE BE 00 BD BD BD 00 BC BC BC 00 BB BB BB 00
BA BA BA 00 B9 B9 B9 00 B8 B8 B8 00 B7 B7 B7 00
B6 B6 B6 00 B5 B5 B5 00 B4 B4 B4 00 B3 B3 B3 00
B2 B2 B2 00 B1 B1 B1 00 B0 B0 B0 00 AF AF AF 00
AE AE AE 00 AD AD AD 00 AC AC AC 00 AB AB AB 00
AA AA AA 00 A9 A9 A9 00 A8 A8 A8 00 A7 A7 A7 00
A6 A6 A6 00 A5 A5 A5 00 A4 A4 A4 00 A3 A3 A3 00
A2 A2 A2 00 A1 A1 A1 00 A0 A0 A0 00 9F 9F 9F 00
9E 9E 9E 00 9D 9D 9D 00 9C 9C 9C 00 9B 9B 9B 00
9A 9A 9A 00 99 99 99 00 98 98 98 00 97 97 97 00
96 96 96 00 95 95 95 00 94 94 94 00 93 93 93 00
92 92 92 00 91 91 91 00 90 90 90 00 8F 8F 8F 00
8E 8E 8E 00 8D 8D 8D 00 8C 8C 8C 00 8B 8B 8B 00
8A 8A 8A 00 89 89 89 00 88 88 88 00 87 87 87 00
86 86 86 00 85 85 85 00 84 84 84 00 83 83 83 00
82 82 82 00 81 81 81 00 80 80 80 00 7F 7F 7F 00
7E 7E 7E 00 7D 7D 7D 00 7C 7C 7C 00 7B 7B 7B 00
7A 7A 7A 00 79 79 79 00 78 78 78 00 77 77 77 00
76 76 76 00 75 75 75 00 74 74 74 00 73 73 73 00
72 72 72 00 71 71 71 00 70 70 70 00 6F 6F 6F 00
6E 6E 6E 00 6D 6D 6D 00 6C 6C 6C 00 6B 6B 6B 00
6A 6A 6A 00 69 69 69 00 68 68 68 00 67 67 67 00
66 66 66 00 65 65 65 00 64 64 64 00 63 63 63 00
62 62 62 00 61 61 61 00 60 60 60 00 5F 5F 5F 00
5E 5E 5E 00 5D 5D 5D 00 5C 5C 5C 00 5B 5B 5B 00
5A 5A 5A 00 59 59 59 00 58 58 58 00 57 57 57 00
56 56 56 00 55 55 55 00 54 54 54 00 53 53 53 00
52 52 52 00 51 51 51 00 50 50 50 00 4F 4F 4F 00
4E 4E 4E 00 4D 4D 4D 00 4C 4C 4C 00 4B 4B 4B 00
4A 4A 4A 00 49 49 49 00 48 48 48 00 47 47 47 00
46 46 46 00 45 45 45 00 44 44 44 00 43 43 43 00
42 42 42 00 41 41 41 00 40 40 40 00 3F 3F 3F 00
3E 3E 3E 00 3D 3D 3D 00 3C 3C 3C 00 3B 3B 3B 00
3A 3A 3A 00 39 39 39 00 38 38 38 00 37 37 37 00
36 36 36 00 35 35 35 00 34 34 34 00 33 33 33 00
32 32 32 00 31 31 31 00 30 30 30 00 2F 2F 2F 00
2E 2E 2E 00 2D 2D 2D 00 2C 2C 2C 00 2B 2B 2B 00
2A 2A 2A 00 29 29 29 00 28 28 28 00 27 27 27 00
26 26 26 00 25 25 25 00 24 24 24 00 23 23 23 00
22 22 22 00 21 21 21 00 20 20 20 00 1F 1F 1F 00
1E 1E 1E 00 1D 1D 1D 00 1C 1C 1C 00 1B 1B 1B 00
1A 1A 1A 00 19 19 19 00 18 18 18 00 17 17 17 00
16 16 16 00 15 15 15 00 14 14 14 00 13 13 13 00
12 12 12 00 11 11 11 00 10 10 10 00 0F 0F 0F 00
0E 0E 0E 00 0D 0D 0D 00 0C 0C 0C 00 0B 0B 0B 00
0A 0A 0A 00 09 09 09 00 08 08 08 00 07 07 07 00
06 06 06 00 05 05 05 00 04 04 04 00 03 03 03 00
02 02 02 00 01 01 01 00 00 00 00 00 00 42 9D 00
00 43 9D 00 01 44 9E 00 01 44 9E 00 02 45 9F 00
02 46 9F 00 02 47 A0 00 03 48 A0 00 03 48 A1 00
04 49 A1 00 04 4A A1 00 04 4B A2 00 05 4C A2 00
05 4C A3 00 05 4D A3 00 06 4E A4 00 06 4F A4 00
07 4F A4 00 07 50 A5 00 07 51 A5 00 08 52 A6 00
08 53 A6 00 09 53 A7 00 09 54 A7 00 09 55 A8 00
0A 56 A8 00 0A 57 A8 00 0B 57 A9 00 0B 58 A9 00
0B 59 AA 00 0C 5A AA 00 0C 5B AB 00 0D 5B AB 00
0D 5C AB 00 0D 5D AC 00 0E 5E AC 00 0E 5F AD 00
0E 5F AD 00 0F 60 AE 00 0F 61 AE 00 10 62 AF 00
10 63 AF 00 10 63 AF 00 11 64 B0 00 11 65 B0 00
12 66 B1 00 12 66 B1 00 12 67 B2 00 13 68 B2 00
13 69 B2 00 14 6A B3 00 14 6A B3 00 14 6B B4 00
15 6C B4 00 15 6D B5 00 16 6E B5 00 16 6E B6 00
16 6F B6 00 17 70 B6 00 17 71 B7 00 17 72 B7 00
18 72 B8 00 18 73 B8 00 19 74 B9 00 19 75 B9 00
19 76 BA 00 1A 76 BA 00 1A 77 BA 00 1B 78 BB 00
1B 79 BB 00 1B 79 BC 00 1C 7A BC 00 1C 7B BD 00
1D 7C BD 00 1D 7D BD 00 1D 7D BE 00 1E 7E BE 00
1E 7F BF 00 1F 80 BF 00 1F 81 C0 00 1F 81 C0 00
20 82 C1 00 20 83 C1 00 20 84 C1 00 21 85 C2 00
21 86 C2 00 22 86 C3 00 22 87 C3 00 22 88 C4 00
23 89 C4 00 23 8A C5 00 24 8A C5 00 24 8B C5 00
24 8C C6 00 25 8D C6 00 25 8E C7 00 26 8E C7 00
26 8F C8 00 26 90 C8 00 27 91 C9 00 27 92 C9 00
28 92 C9 00 28 93 CA 00 28 94 CA 00 29 95 CB 00
29 96 CB 00 2A 96 CC 00 2A 97 CC 00 2A 98 CD 00
2B 99 CD 00 2B 9A CD 00 2C 9A CE 00 2C 9B CE 00
2C 9C CF 00 2D 9D CF 00 2D 9E D0 00 2E 9F D0 00
2E 9F D1 00 2E A0 D1 00 2F A1 D2 00 2F A2 D2 00
30 A3 D2 00 30 A3 D3 00 30 A4 D3 00 31 A5 D4 00
31 A6 D4 00 32 A7 D5 00 32 A7 D5 00 32 A8 D6 00
33 A9 D6 00 33 AA D7 00 34 AB D7 00 34 AC D7 00
34 AC D8 00 35 AD D8 00 35 AE D9 00 36 AF D9 00
36 B0 DA 00 37 B1 DA 00 37 B1 DB 00 37 B2 DB 00
38 B3 DC 00 38 B4 DC 00 39 B5 DC 00 39 B6 DD 00
39 B6 DD 00 3A B7 DE 00 3A B8 DE 00 3B B9 DF 00
3B BA DF 00 3B BA E0 00 3C BB E0 00 3C BC E1 00
3D BD E1 00 3D BE E1 00 3D BF E2 00 3E BF E2 00
3E C0 E3 00 3F C1 E3 00 3F C2 E4 00 40 C3 E4 00
40 C4 E5 00 40 C4 E5 00 41 C5 E6 00 41 C6 E6 00
42 C7 E7 00 42 C8 E7 00 42 C9 E7 00 43 C9 E8 00
43 CA E8 00 44 CB E9 00 44 CC E9 00 44 CD EA 00
45 CE EA 00 45 CF EB 00 46 CF EB 00 46 D0 EC 00
47 D1 EC 00 47 D2 ED 00 47 D3 ED 00 48 D4 EE 00
48 D4 EE 00 49 D5 EE 00 49 D6 EF 00 49 D7 EF 00
4A D8 F0 00 4A D9 F0 00 4B D9 F1 00 4B DA F1 00
4C DB F2 00 4C DC F2 00 4C DD F3 00 4D DE F3 00
4D DF F4 00 4E DF F4 00 4E E0 F5 00 4E E1 F5 00
4F E2 F5 00 4F E3 F6 00 50 E4 F6 00 50 E5 F7 00
51 E5 F7 00 51 E6 F8 00 51 E7 F8 00 52 E8 F9 00
52 E9 F9 00 53 EA FA 00 53 EB FA 00 54 EB FB 00
54 EC FB 00 54 ED FC 00 55 EE FC 00 55 EF FD 00
56 F0 FD 00 56 F0 FE 00 56 F1 FE 00 57 F2 FE 00
57 F3 FF 00 5C F4 FF 00 62 F4 FF 00 68 F4 FF 00
6D F5 FF 00 72 F5 FF 00 77 F6 FF 00 7C F6 FF 00
80 F6 FF 00 85 F7 FF 00 89 F7 FF 00 8E F8 FF 00
92 F8 FF 00 96 F8 FF 00 9B F9 FF 00 9F F9 FF 00
A2 F9 FF 00 A7 FA FF 00 AA FA FF 00 AE FA FF 00
B2 FA FF 00 B6 FB FF 00 B9 FB FF 00 BD FB FF 00
C1 FC FF 00 C4 FC FF 00 C7 FC FF 00 CB FC FF 00
CE FD FF 00 D2 FD FF 00 D5 FD FF 00 D8 FD FF 00
DB FE FF 00 DE FE FF 00 E2 FE FF 00 E5 FF FF 00
E8 FF FF 00 EB FF FF 00 EE FF FF 00 FC 8D 59 00
FC 8E 5A 00 FC 8F 5B 00 FC 90 5B 00 FC 91 5C 00
FC 91 5D 00 FC 92 5E 00 FC 93 5F 00 FC 94 5F 00
FC 95 60 00 FC 96 61 00 FC 97 62 00 FC 98 63 00
FC 99 63 00 FC 9A 64 00 FC 9A 65 00 FC 9B 66 00
FC 9C 67 00 FC 9D 67 00 FC 9E 68 00 FC 9F 69 00
FC A0 6A 00 FD A1 6B 00 FD A2 6B 00 FD A2 6C 00
FD A3 6D 00 FD A4 6E 00 FD A5 6F 00 FD A6 6F 00
FD A7 70 00 FD A8 71 00 FD A9 72 00 FD AA 73 00
FD AB 73 00 FD AB 74 00 FD AC 75 00 FD AD 76 00
FD AE 77 00 FD AF 77 00 FD B0 78 00 FD B1 79 00
FD B2 7A 00 FD B3 7B 00 FD B3 7B 00 FD B4 7C 00
FD B5 7D 00 FD B6 7E 00 FD B7 7F 00 FD B8 7F 00
FD B9 80 00 FD BA 81 00 FD BB 82 00 FD BB 83 00
FD BC 83 00 FD BD 84 00 FD BE 85 00 FD BF 86 00
FD C0 87 00 FD C1 87 00 FD C2 88 00 FD C3 89 00
FD C4 8A 00 FD C4 8B 00 FD C5 8B 00 FE C6 8C 00
FE C7 8D 00 FE C8 8E 00 FE C9 8F 00 FE CA 8F 00
FE CB 90 00 FE CC 91 00 FE CC 92 00 FE CD 93 00
FE CE 93 00 FE CF 94 00 FE D0 95 00 FE D1 96 00
FE D2 97 00 FE D3 97 00 FE D4 98 00 FE D5 99 00
FE D5 9A 00 FE D6 9B 00 FE D7 9B 00 FE D8 9C 00
FE D9 9D 00 FE DA 9E 00 FE DB 9F 00 FE DC 9F 00
FE DD A0 00 FE DD A1 00 FE DE A2 00 FE DF A3 00
FE E0 A3 00 FE E1 A4 00 FE E2 A5 00 FE E3 A6 00
FE E4 A7 00 FE E5 A7 00 FE E6 A8 00 FE E6 A9 00
FE E7 AA 00 FE E8 AB 00 FE E9 AB 00 FE EA AC 00
FE EB AD 00 FE EC AE 00 FF ED AF 00 FF EE AF 00
FF EE B0 00 FF EF B1 00 FF F0 B2 00 FF F1 B3 00
FF F2 B3 00 FF F3 B4 00 FF F4 B5 00 FF F5 B6 00
FF F6 B7 00 FF F7 B7 00 FF F7 B8 00 FF F8 B9 00
FF F9 BA 00 FF FA BB 00 FF FB BB 00 FF FC BC 00
FF FD BD 00 FF FE BE 00 FF FF BF 00 FF FF BF 00
FE FF BE 00 FD FE BE 00 FC FE BE 00 FB FE BD 00
FB FD BD 00 FA FD BD 00 F9 FD BC 00 F8 FC BC 00
F7 FC BC 00 F7 FC BB 00 F6 FB BB 00 F5 FB BB 00
F4 FB BA 00 F3 FA BA 00 F3 FA BA 00 F2 FA B9 00
F1 F9 B9 00 F0 F9 B9 00 EF F9 B8 00 EF F8 B8 00
EE F8 B8 00 ED F8 B7 00 EC F7 B7 00 EB F7 B7 00
EB F7 B6 00 EA F6 B6 00 E9 F6 B6 00 E8 F6 B5 00
E7 F5 B5 00 E7 F5 B5 00 E6 F5 B4 00 E5 F4 B4 00
E4 F4 B4 00 E3 F4 B3 00 E3 F3 B3 00 E2 F3 B3 00
E1 F3 B2 00 E0 F2 B2 00 DF F2 B2 00 DF F2 B1 00
DE F1 B1 00 DD F1 B1 00 DC F1 B0 00 DB F0 B0 00
DB F0 B0 00 DA F0 AF 00 D9 EF AF 00 D8 EF AF 00
D7 EF AE 00 D7 EE AE 00 D6 EE AE 00 D5 EE AD 00
D4 ED AD 00 D3 ED AD 00 D3 ED AC 00 D2 EC AC 00
D1 EC AC 00 D0 EC AB 00 CF EB AB 00 CF EB AB 00
CE EB AA 00 CD EA AA 00 CC EA AA 00 CB EA A9 00
CB E9 A9 00 CA E9 A9 00 C9 E9 A8 00 C8 E8 A8 00
C7 E8 A8 00 C7 E8 A7 00 C6 E7 A7 00 C5 E7 A7 00
C4 E7 A6 00 C3 E6 A6 00 C3 E6 A6 00 C2 E6 A5 00
C1 E5 A5 00 C0 E5 A5 00 BF E5 A4 00 BF E4 A4 00
BE E4 A4 00 BD E4 A3 00 BC E3 A3 00 BB E3 A3 00
BB E3 A2 00 BA E3 A2 00 B9 E2 A1 00 B8 E2 A1 00
B7 E2 A1 00 B7 E1 A0 00 B6 E1 A0 00 B5 E1 A0 00
B4 E0 9F 00 B3 E0 9F 00 B3 E0 9F 00 B2 DF 9E 00
B1 DF 9E 00 B0 DF 9E 00 AF DE 9D 00 AF DE 9D 00
AE DE 9D 00 AD DD 9C 00 AC DD 9C 00 AB DD 9C 00
AB DC 9B 00 AA DC 9B 00 A9 DC 9B 00 A8 DB 9A 00
A7 DB 9A 00 A7 DB 9A 00 A6 DA 99 00 A5 DA 99 00
A4 DA 99 00 A3 D9 98 00 A3 D9 98 00 A2 D9 98 00
A1 D8 97 00 A0 D8 97 00 9F D8 97 00 9F D7 96 00
9E D7 96 00 9D D7 96 00 9C D6 95 00 9B D6 95 00
9B D6 95 00 9A D5 94 00 99 D5 94 00 FF FF CC 00
FE FE CC 00 FC FE CB 00 FB FD CB 00 F9 FD CA 00
F8 FC CA 00 F6 FC CA 00 F5 FB C9 00 F3 FA C9 00
F2 FA C9 00 F0 F9 C8 00 EF F9 C8 00 ED F8 C7 00
EC F7 C7 00 EA F7 C7 00 E9 F6 C6 00 E7 F6 C6 00
E6 F5 C6 00 E4 F5 C5 00 E3 F4 C5 00 E2 F3 C4 00
E0 F3 C4 00 DF F2 C4 00 DD F2 C3 00 DC F1 C3 00
DA F0 C3 00 D9 F0 C2 00 D7 EF C2 00 D6 EF C1 00
D4 EE C1 00 D3 EE C1 00 D1 ED C0 00 D0 EC C0 00
CE EC C0 00 CD EB BF 00 CB EB BF 00 CA EA BE 00
C8 EA BE 00 C7 E9 BE 00 C5 E8 BD 00 C4 E8 BD 00
C3 E7 BD 00 C1 E7 BC 00 C0 E6 BC 00 BE E5 BB 00
BD E5 BB 00 BB E4 BB 00 BA E4 BA 00 B8 E3 BA 00
B7 E3 BA 00 B5 E2 B9 00 B4 E1 B9 00 B2 E1 B8 00
B1 E0 B8 00 AF E0 B8 00 AE DF B7 00 AC DE B7 00
AB DE B7 00 A9 DD B6 00 A8 DD B6 00 A7 DC B5 00
A5 DC B5 00 A4 DB B5 00 A2 DA B4 00 A1 DA B4 00
9F D9 B4 00 9E D9 B5 00 9C D8 B5 00 9B D8 B5 00
99 D7 B5 00 98 D6 B6 00 96 D6 B6 00 95 D5 B6 00
93 D5 B6 00 92 D4 B7 00 90 D4 B7 00 8F D3 B7 00
8D D3 B7 00 8C D2 B8 00 8A D1 B8 00 89 D1 B8 00
87 D0 B8 00 86 D0 B9 00 84 CF B9 00 83 CF B9 00
81 CE B9 00 7F CD BA 00 7E CD BA 00 7C CC BA 00
7B CC BA 00 79 CB BB 00 78 CB BB 00 76 CA BB 00
75 C9 BB 00 73 C9 BC 00 72 C8 BC 00 70 C8 BC 00
6F C7 BC 00 6D C7 BD 00 6C C6 BD 00 6A C6 BD 00
69 C5 BD 00 67 C4 BE 00 66 C4 BE 00 64 C3 BE 00
63 C3 BE 00 61 C2 BF 00 60 C2 BF 00 5E C1 BF 00
5D C0 BF 00 5B C0 C0 00 5A BF C0 00 58 BF C0 00
57 BE C0 00 55 BE C1 00 54 BD C1 00 52 BC C1 00
51 BC C1 00 4F BB C2 00 4E BB C2 00 4C BA C2 00
4B BA C2 00 49 B9 C3 00 48 B9 C3 00 46 B8 C3 00
45 B7 C3 00 43 B7 C4 00 42 B6 C4 00 41 B6 C4 00
41 B5 C4 00 40 B4 C4 00 40 B3 C3 00 40 B2 C3 00
3F B1 C3 00 3F B0 C3 00 3F B0 C3 00 3E AF C2 00
3E AE C2 00 3E AD C2 00 3D AC C2 00 3D AB C2 00
3D AA C1 00 3C A9 C1 00 3C A9 C1 00 3C A8 C1 00
3B A7 C1 00 3B A6 C1 00 3B A5 C0 00 3A A4 C0 00
3A A3 C0 00 3A A3 C0 00 39 A2 C0 00 39 A1 BF 00
39 A0 BF 00 38 9F BF 00 38 9E BF 00 38 9D BF 00
37 9D BE 00 37 9C BE 00 37 9B BE 00 36 9A BE 00
36 99 BE 00 36 98 BE 00 35 97 BD 00 35 97 BD 00
35 96 BD 00 34 95 BD 00 34 94 BD 00 34 93 BC 00
33 92 BC 00 33 91 BC 00 33 90 BC 00 32 90 BC 00
32 8F BB 00 32 8E BB 00 31 8D BB 00 31 8C BB 00
31 8B BB 00 30 8A BA 00 30 8A BA 00 30 89 BA 00
2F 88 BA 00 2F 87 BA 00 2F 86 BA 00 2E 85 B9 00
2E 84 B9 00 2E 84 B9 00 2D 83 B9 00 2D 82 B9 00
2D 81 B8 00 2C 80 B8 00 2C 7F B8 00 2C 7E B8 00
2C 7D B7 00 2C 7C B6 00 2C 7B B6 00 2B 79 B5 00
2B 78 B5 00 2B 77 B4 00 2B 76 B4 00 2B 75 B3 00
2B 74 B2 00 2B 72 B2 00 2B 71 B1 00 2B 70 B1 00
2A 6F B0 00 2A 6E B0 00 2A 6C AF 00 2A 6B AF 00
2A 6A AE 00 2A 69 AD 00 2A 68 AD 00 2A 67 AC 00
2A 65 AC 00 2A 64 AB 00 29 63 AB 00 29 62 AA 00
29 61 A9 00 29 60 A9 00 29 5E A8 00 29 5D A8 00
29 5C A7 00 29 5B A7 00 29 5A A6 00 28 58 A6 00
28 57 A5 00 28 56 A4 00 28 55 A4 00 28 54 A3 00
28 53 A3 00 28 51 A2 00 28 50 A2 00 28 4F A1 00
27 4E A0 00 27 4D A0 00 27 4C 9F 00 27 4A 9F 00
27 49 9E 00 27 48 9E 00 27 47 9D 00 27 46 9C 00
27 44 9C 00 26 43 9B 00 26 42 9B 00 26 41 9A 00
26 40 9A 00 26 3F 99 00 26 3D 99 00 26 3C 98 00
26 3B 97 00 26 3A 97 00 25 39 96 00 25 38 96 00
25 36 95 00 25 35 95 00 25 34 94 00 FE EB E2 00
FE EA E1 00 FE E9 E1 00 FE E8 E0 00 FE E7 DF 00
FE E6 DE 00 FE E5 DE 00 FE E4 DD 00 FE E3 DC 00
FE E2 DB 00 FD E1 DB 00 FD E0 DA 00 FD DF D9 00
FD DE D8 00 FD DD D8 00 FD DC D7 00 FD DB D6 00
FD DA D6 00 FD D9 D5 00 FD D8 D4 00 FD D7 D3 00
FD D6 D3 00 FD D5 D2 00 FD D4 D1 00 FD D3 D0 00
FD D2 D0 00 FD D1 CF 00 FD D0 CE 00 FD D0 CE 00
FC CE CD 00 FC CD CC 00 FC CC CB 00 FC CB CA 00
FC CB CA 00 FC C9 C9 00 FC C8 C8 00 FC C7 C8 00
FC C6 C7 00 FC C5 C6 00 FC C4 C5 00 FC C3 C4 00
FC C2 C4 00 FC C1 C3 00 FC C0 C2 00 FC BF C1 00
FC BE C1 00 FC BD C0 00 FB BC BF 00 FB BB BE 00
FB BA BE 00 FB B9 BD 00 FB B8 BC 00 FB B7 BB 00
FB B6 BB 00 FB B5 BA 00 FB B4 B9 00 FB B3 B9 00
FB B2 B8 00 FB B1 B8 00 FB B0 B8 00 FB AF B7 00
FB AE B7 00 FB AD B7 00 FB AB B6 00 FA AA B6 00
FA A9 B6 00 FA A8 B5 00 FA A7 B5 00 FA A6 B5 00
FA A5 B4 00 FA A4 B4 00 FA A3 B3 00 FA A1 B3 00
FA A0 B3 00 FA 9F B2 00 FA 9E B2 00 FA 9D B2 00
FA 9C B1 00 FA 9B B1 00 FA 9A B1 00 FA 98 B0 00
F9 97 B0 00 F9 96 B0 00 F9 95 AF 00 F9 94 AF 00
F9 93 AE 00 F9 91 AE 00 F9 90 AE 00 F9 8F AD 00
F9 8E AD 00 F9 8D AD 00 F9 8B AC 00 F9 8A AC 00
F9 89 AB 00 F9 88 AB 00 F9 87 AB 00 F9 85 AA 00
F8 84 AA 00 F8 83 AA 00 F8 82 A9 00 F8 80 A9 00
F8 7F A8 00 F8 7E A8 00 F8 7D A8 00 F8 7B A7 00
F8 7A A7 00 F8 79 A6 00 F8 78 A6 00 F8 76 A6 00
F8 75 A5 00 F8 74 A5 00 F8 72 A4 00 F7 71 A4 00
F7 70 A3 00 F7 6E A3 00 F7 6D A3 00 F7 6B A2 00
F7 6A A2 00 F7 69 A1 00 F7 67 A1 00 F6 66 A1 00
F5 66 A0 00 F5 65 A0 00 F4 64 A0 00 F4 63 9F 00
F3 62 9F 00 F2 61 9F 00 F2 60 9F 00 F1 5F 9E 00
F0 5E 9E 00 F0 5D 9E 00 EF 5C 9D 00 EE 5B 9D 00
EE 5A 9D 00 ED 59 9C 00 ED 58 9C 00 EC 57 9C 00
EB 56 9C 00 EB 55 9B 00 EA 54 9B 00 E9 53 9B 00
E9 52 9A 00 E8 51 9A 00 E7 50 9A 00 E7 4F 9A 00
E6 4E 99 00 E5 4D 99 00 E5 4C 99 00 E4 4B 98 00
E3 4A 98 00 E3 49 98 00 E2 48 97 00 E1 47 97 00
E1 46 97 00 E0 45 96 00 DF 44 96 00 DF 42 96 00
DE 41 95 00 DD 40 95 00 DD 3F 95 00 DC 3E 95 00
DB 3D 94 00 DA 3C 94 00 DA 3B 94 00 D9 3A 93 00
D8 39 93 00 D8 38 93 00 D7 37 92 00 D6 35 92 00
D5 34 92 00 D5 33 91 00 D4 32 91 00 D3 31 91 00
D3 30 90 00 D2 2F 90 00 D1 2E 90 00 D0 2C 8F 00
D0 2B 8F 00 CF 2A 8E 00 CE 29 8E 00 CD 28 8E 00
CC 26 8D 00 CC 25 8D 00 CB 24 8D 00 CA 23 8C 00
C9 22 8C 00 C8 20 8C 00 C8 1F 8B 00 C7 1E 8B 00
C6 1C 8A 00 C5 1B 8A 00 C4 1B 8A 00 C3 1A 89 00
C2 1A 89 00 C1 19 89 00 BF 19 89 00 BE 19 88 00
BD 18 88 00 BC 18 88 00 BB 17 87 00 BA 17 87 00
B8 17 87 00 B7 16 86 00 B6 16 86 00 B5 15 86 00
B4 15 86 00 B3 15 85 00 B1 14 85 00 B0 14 85 00
AF 13 84 00 AE 13 84 00 AD 13 84 00 AC 12 84 00
AA 12 83 00 A9 11 83 00 A8 11 83 00 A7 11 82 00
A6 10 82 00 A5 10 82 00 A3 0F 81 00 A2 0F 81 00
A1 0F 81 00 A0 0E 81 00 9F 0E 80 00 9E 0D 80 00
9C 0D 80 00 9B 0D 7F 00 9A 0C 7F 00 99 0C 7F 00
98 0B 7F 00 97 0B 7E 00 95 0B 7E 00 94 0A 7E 00
93 0A 7D 00 92 09 7D 00 91 09 7D 00 90 09 7C 00
8F 08 7C 00 8D 08 7C 00 8C 07 7C 00 8B 07 7B 00
8A 07 7B 00 89 06 7B 00 88 06 7A 00 86 05 7A 00
85 05 7A 00 84 05 7A 00 83 04 79 00 82 04 79 00
81 03 79 00 80 03 78 00 7E 03 78 00 7D 02 78 00
7C 02 78 00 7B 01 77 00 7A 01 77 00 0D 08 87 00
11 08 88 00 15 08 89 00 18 08 8A 00 1B 08 8A 00
1E 08 8B 00 21 08 8C 00 24 08 8C 00 26 08 8D 00
29 08 8E 00 2B 08 8E 00 2E 08 8F 00 30 08 8F 00
32 08 90 00 35 08 90 00 37 08 91 00 39 08 91 00
3B 08 92 00 3D 08 92 00 3F 08 93 00 41 08 93 00
43 08 94 00 45 08 94 00 47 08 95 00 49 08 95 00
4B 08 96 00 4D 09 96 00 4F 09 97 00 51 09 97 00
53 09 98 00 54 09 98 00 56 09 98 00 58 09 99 00
5A 09 99 00 5C 09 9A 00 5D 09 9A 00 5F 09 9B 00
61 09 9B 00 63 09 9B 00 64 09 9C 00 66 09 9C 00
68 09 9D 00 69 09 9D 00 6B 09 9D 00 6D 09 9E 00
6F 09 9E 00 70 09 9F 00 72 09 9F 00 74 09 9F 00
75 09 A0 00 77 09 A0 00 79 09 A1 00 7A 09 A1 00
7C 09 A1 00 7E 09 A2 00 7F 09 A2 00 81 09 A3 00
82 09 A3 00 84 09 A3 00 86 09 A4 00 87 09 A4 00
89 09 A5 00 8B 09 A5 00 8C 0A A4 00 8E 0C A3 00
90 0E A1 00 92 10 A0 00 93 12 9F 00 95 13 9D 00
97 15 9C 00 98 17 9B 00 9A 18 9A 00 9B 1A 99 00
9C 1B 98 00 9E 1D 97 00 9F 1E 96 00 A1 1F 95 00
A2 21 93 00 A3 22 92 00 A5 23 92 00 A6 25 91 00
A7 26 90 00 A8 27 8F 00 AA 29 8E 00 AB 2A 8D 00
AC 2B 8C 00 AD 2C 8B 00 AE 2E 8A 00 AF 2F 89 00
B1 30 88 00 B2 31 87 00 B3 32 87 00 B4 34 86 00
B5 35 85 00 B6 36 84 00 B7 37 83 00 B8 38 82 00
BA 39 81 00 BB 3A 81 00 BC 3C 80 00 BD 3D 7F 00
BE 3E 7E 00 BF 3F 7D 00 C0 40 7D 00 C1 41 7C 00
C2 42 7B 00 C3 43 7A 00 C4 44 79 00 C5 45 79 00
C6 46 78 00 C7 47 77 00 C8 49 76 00 C9 4A 76 00
CA 4B 75 00 CB 4C 74 00 CC 4D 73 00 CD 4E 72 00
CE 4F 72 00 CF 50 71 00 D0 51 70 00 D1 52 6F 00
D2 53 6F 00 D3 54 6E 00 D4 55 6D 00 D5 56 6D 00
D6 57 6C 00 D7 58 6B 00 D8 59 6A 00 D9 5A 6A 00
DA 5B 69 00 DB 5C 68 00 DB 5D 67 00 DC 5F 66 00
DD 60 65 00 DD 61 65 00 DE 63 64 00 DE 64 63 00
DF 65 62 00 DF 67 61 00 E0 68 60 00 E0 69 60 00
E1 6B 5F 00 E1 6C 5E 00 E2 6D 5D 00 E2 6F 5C 00
E2 70 5C 00 E3 71 5B 00 E3 73 5A 00 E4 74 59 00
E4 75 58 00 E5 76 58 00 E5 78 57 00 E6 79 56 00
E6 7A 55 00 E7 7B 54 00 E7 7D 54 00 E8 7E 53 00
E8 7F 52 00 E9 80 51 00 E9 81 51 00 E9 83 50 00
EA 84 4F 00 EA 85 4E 00 EB 86 4E 00 EB 88 4D 00
EC 89 4C 00 EC 8A 4B 00 ED 8B 4B 00 ED 8C 4A 00
EE 8D 49 00 EE 8F 48 00 EE 90 48 00 EF 91 47 00
EF 92 46 00 F0 93 45 00 F0 95 45 00 F1 96 44 00
F1 97 43 00 F2 98 42 00 F2 99 42 00 F2 9A 41 00
F3 9C 40 00 F3 9D 40 00 F4 9E 3F 00 F4 9F 3E 00
F5 A0 3D 00 F5 A1 3D 00 F5 A2 3C 00 F6 A4 3B 00
F6 A5 3B 00 F7 A6 3A 00 F7 A7 39 00 F8 A8 38 00
F8 A9 38 00 F8 AA 37 00 F9 AC 36 00 F9 AD 36 00
FA AE 35 00 FA AF 34 00 FB B0 33 00 FB B1 33 00
FB B2 32 00 FC B4 31 00 FC B5 31 00 FD B6 30 00
FD B7 2F 00 FE B8 2E 00 FE B9 2E 00 FE BA 2D 00
FF BB 2C 00 FF BD 2C 00 FE BE 2C 00 FE C0 2B 00
FE C1 2B 00 FD C2 2B 00 FD C4 2B 00 FD C5 2A 00
FC C7 2A 00 FC C8 2A 00 FC C9 2A 00 FB CB 29 00
FB CC 29 00 FB CE 29 00 FA CF 29 00 FA D0 28 00
FA D2 28 00 F9 D3 28 00 F9 D4 28 00 F9 D6 27 00
F8 D7 27 00 F8 D8 27 00 F8 DA 27 00 F7 DB 26 00
F7 DD 26 00 F7 DE 26 00 F6 DF 26 00 F6 E0 25 00
F6 E2 25 00 F5 E3 25 00 F5 E4 25 00 F5 E6 24 00
F4 E7 24 00 F4 E8 24 00 F4 EA 24 00 F3 EB 24 00
F3 EC 23 00 F3 EE 23 00 F3 EF 23 00 F2 F0 23 00
F2 F1 22 00 F2 F3 22 00 F1 F4 22 00 F1 F5 22 00
F1 F6 21 00 F0 F8 21 00 F0 F9 21 00 FF 00 00 00
FF 06 00 00 FF 0C 00 00 FF 12 00 00 FF 18 00 00
FF 1E 00 00 FF 24 00 00 FF 2A 00 00 FF 30 00 00
FF 36 00 00 FF 3C 00 00 FF 42 00 00 FF 48 00 00
FF 4E 00 00 FF 54 00 00 FF 5A 00 00 FF 60 00 00
FF 66 00 00 FF 6C 00 00 FF 72 00 00 FF 78 00 00
FF 7E 00 00 FF 84 00 00 FF 8A 00 00 FF 90 00 00
FF 96 00 00 FF 9C 00 00 FF A2 00 00 FF A8 00 00
FF AE 00 00 FF B4 00 00 FF BA 00 00 FF C0 00 00
FF C6 00 00 FF CC 00 00 FF D2 00 00 FF D8 00 00
FF DE 00 00 FF E4 00 00 FF EA 00 00 FF F0 00 00
FF F6 00 00 FF FC 00 00 FC FF 00 00 F6 FF 00 00
F0 FF 00 00 EA FF 00 00 E4 FF 00 00 DE FF 00 00
D8 FF 00 00 D2 FF 00 00 CC FF 00 00 C6 FF 00 00
C0 FF 00 00 BA FF 00 00 B4 FF 00 00 AE FF 00 00
A8 FF 00 00 A2 FF 00 00 9C FF 00 00 96 FF 00 00
90 FF 00 00 8A FF 00 00 84 FF 00 00 7E FF 00 00
78 FF 00 00 72 FF 00 00 6C FF 00 00 66 FF 00 00
60 FF 00 00 5A FF 00 00 54 FF 00 00 4E FF 00 00
48 FF 00 00 42 FF 00 00 3C FF 00 00 36 FF 00 00
30 FF 00 00 2A FF 00 00 24 FF 00 00 1E FF 00 00
18 FF 00 00 12 FF 00 00 0C FF 00 00 06 FF 00 00
00 FF 00 00 00 FF 06 00 00 FF 0C 00 00 FF 12 00
00 FF 18 00 00 FF 1E 00 00 FF 24 00 00 FF 2A 00
00 FF 30 00 00 FF 36 00 00 FF 3C 00 00 FF 42 00
00 FF 48 00 00 FF 4E 00 00 FF 54 00 00 FF 5A 00
00 FF 60 00 00 FF 66 00 00 FF 6C 00 00 FF 72 00
00 FF 78 00 00 FF 7E 00 00 FF 84 00 00 FF 8A 00
00 FF 90 00 00 FF 96 00 00 FF 9C 00 00 FF A2 00
00 FF A8 00 00 FF AE 00 00 FF B4 00 00 FF BA 00
00 FF C0 00 00 FF C6 00 00 FF CC 00 00 FF D2 00
00 FF D8 00 00 FF DE 00 00 FF E4 00 00 FF EA 00
00 FF F0 00 00 FF F6 00 00 FF FC 00 00 FC FF 00
00 F6 FF 00 00 F0 FF 00 00 EA FF 00 00 E4 FF 00
00 DE FF 00 00 D8 FF 00 00 D2 FF 00 00 CC FF 00
00 C6 FF 00 00 C0 FF 00 00 BA FF 00 00 B4 FF 00
00 AE FF 00 00 A8 FF 00 00 A2 FF 00 00 9C FF 00
00 96 FF 00 00 90 FF 00 00 8A FF 00 00 84 FF 00
00 7E FF 00 00 78 FF 00 00 72 FF 00 00 6C FF 00
00 66 FF 00 00 60 FF 00 00 5A FF 00 00 54 FF 00
00 4E FF 00 00 48 FF 00 00 42 FF 00 00 3C FF 00
00 36 FF 00 00 30 FF 00 00 2A FF 00 00 24 FF 00
00 1E FF 00 00 18 FF 00 00 12 FF 00 00 0C FF 00
00 06 FF 00 00 00 FF 00 06 00 FF 00 0C 00 FF 00
12 00 FF 00 18 00 FF 00 1E 00 FF 00 24 00 FF 00
2A 00 FF 00 30 00 FF 00 36 00 FF 00 3C 00 FF 00
42 00 FF 00 48 00 FF 00 4E 00 FF 00 54 00 FF 00
5A 00 FF 00 60 00 FF 00 66 00 FF 00 6C 00 FF 00
72 00 FF 00 78 00 FF 00 7E 00 FF 00 84 00 FF 00
8A 00 FF 00 90 00 FF 00 96 00 FF 00 9C 00 FF 00
A2 00 FF 00 A8 00 FF 00 AE 00 FF 00 B4 00 FF 00
BA 00 FF 00 C0 00 FF 00 C6 00 FF 00 CC 00 FF 00
D2 00 FF 00 D8 00 FF 00 DE 00 FF 00 E4 00 FF 00
EA 00 FF 00 F0 00 FF 00 F6 00 FF 00 FC 00 FF 00
FF 00 FC 00 FF 00 F6 00 FF 00 F0 00 FF 00 EA 00
FF 00 E4 00 FF 00 DE 00 FF 00 D8 00 FF 00 D2 00
FF 00 CC 00 FF 00 C6 00 FF 00 C0 00 FF 00 BA 00
FF 00 B4 00 FF 00 AE 00 FF 00 A8 00 FF 00 A2 00
FF 00 9C 00 FF 00 96 00 FF 00 90 00 FF 00 8A 00
FF 00 84 00 FE 00 7F 00 FE 00 79 00 FE 00 73 00
FE 00 6D 00 FE 00 67 00 FE 00 61 00 FE 00 5B 00
FE 00 55 00 FE 00 4F 00 FE 00 49 00 FE 00 43 00
FE 00 3D 00 FE 00 37 00 FE 00 31 00 FE 00 2B 00
FE 00 25 00 FE 00 1F 00 FE 00 19 00 FE 00 13 00
FE 00 0D 00 FE 00 07 00 FE 00 01 00
@00002C5C
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
84 D3 FF FF 18 00 00 00 00 00 00 00
@00002C88
04 00 01 80 00 00 00 80 9A 99 A3 FC 9A 99 03 FA
