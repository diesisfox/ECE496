/**** write_top_decl_start_and_interfaces output below ****/

module top(
    input clock, reset_n,
    output cpu_trap,
    input logic CLOCK_50,
    output logic [7:0]VGA_R,
    output logic [7:0]VGA_G,
    output logic [7:0]VGA_B,
    output logic VGA_CLK,
    output logic VGA_SYNC_N,
    output logic VGA_BLANK_N,
    output logic VGA_HS,
    output logic VGA_VS,
    input logic [9:0]SW,
    input logic [3:0]KEY,
    output logic [9:0]LEDR,
    inout logic GPIO_0[0],
    inout logic GPIO_0[1],
    inout logic GPIO_0[2],
    inout logic GPIO_0[3],
    inout logic GPIO_0[4],
    inout logic GPIO_0[5],
    inout logic GPIO_0[6]
);

AXI5_Lite_IF M_IF ();

Simple_Worker_Mem_IF mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_if0();

Simple_Worker_Mem_IF IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if0();

IP_VGA_IF IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1();
tran(CLOCK_50, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.CLOCK_50);
tran([7:0]VGA_R, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_R);
tran([7:0]VGA_G, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_G);
tran([7:0]VGA_B, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_B);
tran(VGA_CLK, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_CLK);
tran(VGA_SYNC_N, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_SYNC_N);
tran(VGA_BLANK_N, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_BLANK_N);
tran(VGA_HS, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_HS);
tran(VGA_VS, IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1.VGA_VS);

Simple_Worker_Mem_IF IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if0();

IP_GPIO_IF IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if1();
tran([9:0]SW, IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if1.pins);

Simple_Worker_Mem_IF IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if0();

IP_GPIO_IF IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if1();
tran([3:0]KEY, IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if1.pins);

Simple_Worker_Mem_IF IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if0();

IP_GPIO_IF IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if1();
tran([9:0]LEDR, IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if1.pins);

Simple_Worker_Mem_IF IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if0();

IP_GPIO_IF IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1();
tran(GPIO_0[0], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[0]);
tran(GPIO_0[1], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[1]);
tran(GPIO_0[2], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[2]);
tran(GPIO_0[3], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[3]);
tran(GPIO_0[4], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[4]);
tran(GPIO_0[5], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[5]);
tran(GPIO_0[6], IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1.pins[6]);


/**** write_module_instantiations output below ****/


picorv32_axi #(
    .PROGADDR_RESET(32'h0000_0000),
    .STACKADDR(32'h0000_8000),
    .ENABLE_FAST_MUL(1),
    .ENABLE_DIV(1)
) picorv32_axi_7CB48A78B25546A8AC109ED58AE32A4A (
    .clk(clock),
    .resetn(reset_n),
    .trap(cpu_trap),
    .AXI_IF(M_IF)
);

mem_m10k #(
    .ADDR(32'h0000_0000),
    .N_ADDR_BITS(16),
    .MIF_FILENAME("resources/mandel.mif")
) mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7 (
    .mem_if(mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_if0)
);

IP_VGA_Main #(
    .ADDR(32'h8000_0000),
    .DEPTH(8),
    .W_DIV_1280(1),
    .H_DIV_960(1),
    .VRAM_MIF("resources/peripherals/vga/480_1502934674.inkh_59_melloque_waifu2x_art_scale_tta_1 copy_waifu2x_art_noise3_scale_tta_1 copy 2.png.p256.png.mif"),
    .PALETTE_MIF("resources/peripherals/vga/480_1502934674.inkh_59_melloque_waifu2x_art_scale_tta_1 copy_waifu2x_art_noise3_scale_tta_1 copy 2.png.palette.png.mif")
) IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F (
    .Bus(IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if0),
    .VGA_IF(IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if1)
);

IP_GPIO_Main #(
    .ADDR(32'h8000_0020),
    .PINS(10)
) IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B (
    .Bus(IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if0),
    .Pins(IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if1)
);

IP_GPIO_Main #(
    .ADDR(32'h8000_0030),
    .PINS(4)
) IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689 (
    .Bus(IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if0),
    .Pins(IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if1)
);

IP_GPIO_Main #(
    .ADDR(32'h8000_0040),
    .PINS(10)
) IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D (
    .Bus(IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if0),
    .Pins(IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if1)
);

IP_GPIO_Main #(
    .ADDR(32'h8000_0050),
    .PINS(7)
) IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E (
    .Bus(IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if0),
    .Pins(IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if1)
);


/**** write_controller_and_interconnect_inst output below ****/

    AXI_Controller_Worker mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_controller (
        .AXI_IF(mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_AXI_if0),
        .USER_IF(mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_if0)
    );

    AXI_Controller_Worker IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_controller (
        .AXI_IF(IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_AXI_if0),
        .USER_IF(IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_if0)
    );

    AXI_Controller_Worker IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_controller (
        .AXI_IF(IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_AXI_if0),
        .USER_IF(IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_if0)
    );

    AXI_Controller_Worker IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_controller (
        .AXI_IF(IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_AXI_if0),
        .USER_IF(IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_if0)
    );

    AXI_Controller_Worker IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_controller (
        .AXI_IF(IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_AXI_if0),
        .USER_IF(IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_if0)
    );

    AXI_Controller_Worker IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_controller (
        .AXI_IF(IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_AXI_if0),
        .USER_IF(IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_if0)
    );

    AXI_Interconnect #(
        .mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_base_addr(32'h0000_0000),
        .mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits(16),
        .IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_base_addr(32'h8000_0000),
        .IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits(5),
        .IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_base_addr(32'h8000_0020),
        .IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits(4),
        .IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_base_addr(32'h8000_0030),
        .IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits(4),
        .IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_base_addr(32'h8000_0040),
        .IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits(4),
        .IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_base_addr(32'h8000_0050),
        .IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits(4)
    ) xbar (
        .mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF(mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_AXI_if0),
        .IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF(IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_AXI_if0),
        .IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF(IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_AXI_if0),
        .IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF(IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_AXI_if0),
        .IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF(IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_AXI_if0),
        .IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF(IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_AXI_if0),
        .M_IF(M_IF)
    );


/**** write_top_verilog_end output below ****/


endmodule //top


/**** write_axi_interconnect output below ****/

module AXI_Interconnect #(
    parameter [31:0] mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_base_addr = 32'h0000_0000,
    parameter int mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits = 16,
    parameter [31:0] IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_base_addr = 32'h8000_0000,
    parameter int IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits = 5,
    parameter [31:0] IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_base_addr = 32'h8000_0020,
    parameter int IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits = 4,
    parameter [31:0] IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_base_addr = 32'h8000_0030,
    parameter int IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits = 4,
    parameter [31:0] IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_base_addr = 32'h8000_0040,
    parameter int IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits = 4,
    parameter [31:0] IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_base_addr = 32'h8000_0050,
    parameter int IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits = 4
)(
    AXI5_Lite_IF.WORKER M_IF,
    AXI5_Lite_IF.MANAGER mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF,
    AXI5_Lite_IF.MANAGER IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF,
    AXI5_Lite_IF.MANAGER IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF,
    AXI5_Lite_IF.MANAGER IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF,
    AXI5_Lite_IF.MANAGER IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF,
    AXI5_Lite_IF.MANAGER IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF
);

    // Clock and reset wiring
    assign mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ACLK = M_IF.ACLK;
    assign mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARESETn = M_IF.ARESETn;
    assign IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ACLK = M_IF.ACLK;
    assign IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARESETn = M_IF.ARESETn;
    assign IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ACLK = M_IF.ACLK;
    assign IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARESETn = M_IF.ARESETn;
    assign IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ACLK = M_IF.ACLK;
    assign IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARESETn = M_IF.ARESETn;
    assign IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ACLK = M_IF.ACLK;
    assign IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARESETn = M_IF.ARESETn;
    assign IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ACLK = M_IF.ACLK;
    assign IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARESETn = M_IF.ARESETn;

    logic [31:0] araddr;
    logic [31:0] araddr_latched;
    logic [31:0] araddr_sel;

    logic [31:0] awaddr;
    logic [31:0] awaddr_latched;
    logic [31:0] awaddr_sel;

    assign araddr = M_IF.ARADDR;
    assign awaddr = M_IF.AWADDR;

    enum logic [1:0] {
        READ_IDLE,
        ARADDR_LATCHED,
        AR_DONE
    } read_state;

    // Read state machine
    always_ff @(posedge M_IF.ACLK) begin
        if (M_IF.ARESETn == 1'b0) begin
            read_state <= READ_IDLE;
        end else begin
            case (read_state)
                READ_IDLE : begin
                    if (M_IF.ARREADY && M_IF.ARVALID) begin
                        read_state <= AR_DONE;
                    end else if (M_IF.ARVALID) begin
                        read_state <= ARADDR_LATCHED;
                    end else begin
                        read_state <= READ_IDLE;
                    end
                end
                ARADDR_LATCHED : begin
                    if (M_IF.ARREADY && M_IF.ARVALID) begin
                        read_state <= AR_DONE;
                    end else begin
                        read_state <= ARADDR_LATCHED;
                    end
                end
                AR_DONE : begin
                    if (M_IF.RREADY && M_IF.RVALID) begin
                        read_state <= READ_IDLE;
                    end else begin
                        read_state <= AR_DONE;
                    end
                end
                default : begin
                    read_state <= read_state;
                end
            endcase
        end
    end

    // ARADDR latching
    always_ff @(posedge M_IF.ACLK) begin
        if (M_IF.ARESETn == 1'b0) begin
            araddr_latched <= 32'b0;
        end else begin
            if (M_IF.ARVALID && read_state == READ_IDLE) begin
                araddr_latched <= M_IF.ARADDR;
            end
        end
    end

    // Wiring for araddr_sel, and read XBAR
    always_comb begin
        // Default case - we expect to never hit this
        araddr_sel = 'b0;
        if (read_state == ARADDR_LATCHED || read_state == AR_DONE) begin
            araddr_sel = araddr_latched;
        end else begin
            araddr_sel = araddr;
        end

        // Default tie-offs
        // Manager
        M_IF.ARREADY = 'b0;
        M_IF.RDATA = 'b0;
        M_IF.RRESP = 'b0;
        M_IF.RVALID = 'b0;
        M_IF.RID = 'b0;

        // mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARADDR = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARPROT = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARVALID = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARSIZE = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARID = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RREADY = 'b0;

        // IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARADDR = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARPROT = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARVALID = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARSIZE = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARID = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RREADY = 'b0;

        // IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARADDR = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARPROT = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARVALID = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARSIZE = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARID = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RREADY = 'b0;

        // IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARADDR = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARPROT = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARVALID = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARSIZE = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARID = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RREADY = 'b0;

        // IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARADDR = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARPROT = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARVALID = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARSIZE = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARID = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RREADY = 'b0;

        // IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARADDR = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARPROT = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARVALID = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARSIZE = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARID = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RREADY = 'b0;

        if (araddr_sel[31:mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits] == mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_base_addr[31:mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits]) begin
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARADDR = M_IF.ARADDR;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARPROT = M_IF.ARPROT;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARREADY;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARSIZE = M_IF.ARSIZE;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.ARID = M_IF.ARID;
            M_IF.RDATA = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RDATA;
            M_IF.RRESP = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RRESP;
            M_IF.RVALID = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RVALID;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RREADY = M_IF.RREADY;
            M_IF.RID = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.RID;
        end else if (araddr_sel[31:IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits] == IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_base_addr[31:IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits]) begin
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARADDR = M_IF.ARADDR;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARPROT = M_IF.ARPROT;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARREADY;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARSIZE = M_IF.ARSIZE;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.ARID = M_IF.ARID;
            M_IF.RDATA = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RDATA;
            M_IF.RRESP = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RRESP;
            M_IF.RVALID = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RVALID;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RREADY = M_IF.RREADY;
            M_IF.RID = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.RID;
        end else if (araddr_sel[31:IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits] == IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_base_addr[31:IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits]) begin
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARADDR = M_IF.ARADDR;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARPROT = M_IF.ARPROT;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARREADY;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARSIZE = M_IF.ARSIZE;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.ARID = M_IF.ARID;
            M_IF.RDATA = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RDATA;
            M_IF.RRESP = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RRESP;
            M_IF.RVALID = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RVALID;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RREADY = M_IF.RREADY;
            M_IF.RID = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.RID;
        end else if (araddr_sel[31:IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits] == IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_base_addr[31:IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits]) begin
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARADDR = M_IF.ARADDR;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARPROT = M_IF.ARPROT;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARREADY;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARSIZE = M_IF.ARSIZE;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.ARID = M_IF.ARID;
            M_IF.RDATA = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RDATA;
            M_IF.RRESP = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RRESP;
            M_IF.RVALID = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RVALID;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RREADY = M_IF.RREADY;
            M_IF.RID = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.RID;
        end else if (araddr_sel[31:IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits] == IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_base_addr[31:IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits]) begin
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARADDR = M_IF.ARADDR;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARPROT = M_IF.ARPROT;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARREADY;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARSIZE = M_IF.ARSIZE;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.ARID = M_IF.ARID;
            M_IF.RDATA = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RDATA;
            M_IF.RRESP = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RRESP;
            M_IF.RVALID = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RVALID;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RREADY = M_IF.RREADY;
            M_IF.RID = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.RID;
        end else if (araddr_sel[31:IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits] == IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_base_addr[31:IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits]) begin
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARADDR = M_IF.ARADDR;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARPROT = M_IF.ARPROT;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARVALID = M_IF.ARVALID;
            M_IF.ARREADY = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARREADY;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARSIZE = M_IF.ARSIZE;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.ARID = M_IF.ARID;
            M_IF.RDATA = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RDATA;
            M_IF.RRESP = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RRESP;
            M_IF.RVALID = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RVALID;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RREADY = M_IF.RREADY;
            M_IF.RID = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.RID;
        end
    end

    enum logic [1:0] {
        WRITE_IDLE,
        AWADDR_LATCHED,
        AW_DONE
    } write_state;

    // Write state machine
    always_ff @(posedge M_IF.ACLK) begin
        if (M_IF.ARESETn == 1'b0) begin
            write_state <= WRITE_IDLE;
        end else begin
            case (write_state)
                WRITE_IDLE : begin
                    if (M_IF.AWREADY && M_IF.AWVALID) begin
                        write_state <= AW_DONE;
                    end else if (M_IF.AWVALID) begin
                        write_state <= AWADDR_LATCHED;
                    end else begin
                        write_state <= WRITE_IDLE;
                    end
                end
                AWADDR_LATCHED : begin
                    if (M_IF.AWREADY && M_IF.AWVALID) begin
                        write_state <= AW_DONE;
                    end else begin
                        write_state <= AWADDR_LATCHED;
                    end
                end
                AW_DONE : begin
                    if (M_IF.BREADY && M_IF.BVALID) begin
                        write_state <= WRITE_IDLE;
                    end else begin
                        write_state <= AW_DONE;
                    end
                end
                default : begin
                    write_state <= write_state;
                end
            endcase
        end
    end

    // AWADDR latching
    always_ff @(posedge M_IF.ACLK) begin
        if (M_IF.ARESETn == 1'b0) begin
            awaddr_latched <= 32'b0;
        end else begin
            if (M_IF.AWVALID && write_state == WRITE_IDLE) begin
                awaddr_latched <= awaddr;
            end
        end
    end

    // Wiring for awaddr_sel and write XBAR
    always_comb begin
        awaddr_sel = 'b0;
        if (write_state == AWADDR_LATCHED || write_state == AW_DONE) begin
            awaddr_sel = awaddr_latched;
        end else begin
            awaddr_sel = awaddr;
        end

        // Default tie-offs
        // Manager
        M_IF.AWREADY = 'b0;
        M_IF.WREADY = 'b0;
        M_IF.BRESP = 'b0;
        M_IF.BVALID = 'b0;
        M_IF.BID = 'b0;

        // mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWADDR = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWPROT = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWVALID = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWSIZE = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWID = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WDATA = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WSTRB = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WVALID = 'b0;
        mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.BREADY = 'b0;

        // IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWADDR = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWPROT = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWVALID = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWSIZE = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWID = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WDATA = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WSTRB = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WVALID = 'b0;
        IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.BREADY = 'b0;

        // IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWADDR = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWPROT = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWVALID = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWSIZE = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWID = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WDATA = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WSTRB = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WVALID = 'b0;
        IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.BREADY = 'b0;

        // IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWADDR = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWPROT = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWVALID = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWSIZE = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWID = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WDATA = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WSTRB = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WVALID = 'b0;
        IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.BREADY = 'b0;

        // IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWADDR = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWPROT = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWVALID = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWSIZE = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWID = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WDATA = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WSTRB = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WVALID = 'b0;
        IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.BREADY = 'b0;

        // IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWADDR = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWPROT = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWVALID = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWSIZE = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWID = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WDATA = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WSTRB = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WVALID = 'b0;
        IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.BREADY = 'b0;

        if (awaddr_sel[31:mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits] == mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_base_addr[31:mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_num_bits]) begin
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWADDR = M_IF.AWADDR;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWPROT = M_IF.AWPROT;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWREADY;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWSIZE = M_IF.AWSIZE;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.AWID = M_IF.AWID;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WDATA = M_IF.WDATA;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WSTRB = M_IF.WSTRB;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.WREADY;
            M_IF.BRESP = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.BRESP;
            M_IF.BVALID = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.BVALID;
            mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.BREADY = M_IF.BREADY;
            M_IF.BID = mem_m10k_931897D0B4814B10A0108CB4D8FD8FD7_IF.BID;
        end else if (awaddr_sel[31:IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits] == IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_base_addr[31:IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_num_bits]) begin
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWADDR = M_IF.AWADDR;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWPROT = M_IF.AWPROT;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWREADY;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWSIZE = M_IF.AWSIZE;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.AWID = M_IF.AWID;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WDATA = M_IF.WDATA;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WSTRB = M_IF.WSTRB;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.WREADY;
            M_IF.BRESP = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.BRESP;
            M_IF.BVALID = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.BVALID;
            IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.BREADY = M_IF.BREADY;
            M_IF.BID = IP_VGA_Main_6367E892C4E74E548BDF4DBD747EC45F_IF.BID;
        end else if (awaddr_sel[31:IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits] == IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_base_addr[31:IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_num_bits]) begin
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWADDR = M_IF.AWADDR;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWPROT = M_IF.AWPROT;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWREADY;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWSIZE = M_IF.AWSIZE;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.AWID = M_IF.AWID;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WDATA = M_IF.WDATA;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WSTRB = M_IF.WSTRB;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.WREADY;
            M_IF.BRESP = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.BRESP;
            M_IF.BVALID = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.BVALID;
            IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.BREADY = M_IF.BREADY;
            M_IF.BID = IP_GPIO_Main_EDCBA89957144E9786243CBAB6035F9B_IF.BID;
        end else if (awaddr_sel[31:IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits] == IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_base_addr[31:IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_num_bits]) begin
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWADDR = M_IF.AWADDR;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWPROT = M_IF.AWPROT;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWREADY;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWSIZE = M_IF.AWSIZE;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.AWID = M_IF.AWID;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WDATA = M_IF.WDATA;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WSTRB = M_IF.WSTRB;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.WREADY;
            M_IF.BRESP = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.BRESP;
            M_IF.BVALID = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.BVALID;
            IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.BREADY = M_IF.BREADY;
            M_IF.BID = IP_GPIO_Main_03E7C7957D28435F9FEA43E474E12689_IF.BID;
        end else if (awaddr_sel[31:IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits] == IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_base_addr[31:IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_num_bits]) begin
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWADDR = M_IF.AWADDR;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWPROT = M_IF.AWPROT;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWREADY;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWSIZE = M_IF.AWSIZE;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.AWID = M_IF.AWID;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WDATA = M_IF.WDATA;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WSTRB = M_IF.WSTRB;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.WREADY;
            M_IF.BRESP = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.BRESP;
            M_IF.BVALID = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.BVALID;
            IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.BREADY = M_IF.BREADY;
            M_IF.BID = IP_GPIO_Main_A82B8DF9798D4A83A773B4EB08A2678D_IF.BID;
        end else if (awaddr_sel[31:IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits] == IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_base_addr[31:IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_num_bits]) begin
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWADDR = M_IF.AWADDR;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWPROT = M_IF.AWPROT;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWVALID = M_IF.AWVALID;
            M_IF.AWREADY = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWREADY;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWSIZE = M_IF.AWSIZE;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.AWID = M_IF.AWID;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WDATA = M_IF.WDATA;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WSTRB = M_IF.WSTRB;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WVALID = M_IF.WVALID;
            M_IF.WREADY = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.WREADY;
            M_IF.BRESP = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.BRESP;
            M_IF.BVALID = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.BVALID;
            IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.BREADY = M_IF.BREADY;
            M_IF.BID = IP_GPIO_Main_E55DA6BDF4EC42659239D2DD6B45F15E_IF.BID;
        end
    end

endmodule
