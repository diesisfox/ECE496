module AXI_Controller_Worker ();

endmodule
