@00000000
97 11 00 00 93 81 81 CD 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 80 3D
@00000006
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 A4 FE
23 24 B4 FE 83 25 C4 FE 13 88 05 00 93 D5 F5 41
93 88 05 00 83 25 84 FE 13 86 05 00 93 D5 F5 41
93 86 05 00 33 85 C8 02 B3 85 06 03 B3 05 B5 00
33 05 C8 02 B3 37 C8 02 13 07 05 00 B3 86 F5 00
93 87 06 00 93 96 67 00 13 53 A7 01 33 E3 66 00
93 D3 A7 41 93 07 03 00 13 85 07 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FC 23 2E 11 02
23 2C 81 02 23 2A 91 02 13 04 01 04 23 26 A4 FC
23 24 B4 FC 93 07 F0 FF A3 01 F4 FE A3 07 04 FE
23 24 04 FE 23 22 04 FE 6F 00 C0 07 83 25 84 FE
03 25 84 FE EF F0 DF F4 93 04 05 00 83 25 44 FE
03 25 44 FE EF F0 DF F3 93 07 05 00 B3 87 F4 40
03 27 C4 FC B3 07 F7 00 23 2E F4 FC 83 25 84 FE
37 05 00 08 EF F0 DF F1 93 07 05 00 83 25 44 FE
13 85 07 00 EF F0 DF F0 13 07 05 00 83 27 84 FC
B3 87 E7 00 23 2C F4 FC 83 27 C4 FD 23 24 F4 FE
83 27 84 FD 23 22 F4 FE 83 47 F4 FE 93 87 17 00
A3 07 F4 FE 83 25 84 FE 03 25 84 FE EF F0 5F ED
93 04 05 00 83 25 44 FE 03 25 44 FE EF F0 5F EC
93 07 05 00 33 87 F4 00 B7 07 00 10 63 C8 E7 00
03 47 F4 FE 83 47 34 FE E3 6A F7 F4 83 47 F4 FE
13 85 07 00 83 20 C1 03 03 24 81 03 83 24 41 03
13 01 01 04 67 80 00 00 13 01 01 FC 23 2E 11 02
23 2C 81 02 13 04 01 04 23 26 A4 FC 23 24 B4 FC
23 22 C4 FC 23 20 D4 FC 03 27 84 FC 83 27 C4 FC
33 07 F7 40 B7 A7 01 00 93 85 A7 99 13 05 07 00
EF F0 1F E5 23 2E A4 FC 03 27 C4 FC 83 27 C4 FD
B3 07 F7 00 93 D7 17 40 23 2C F4 FC 03 27 44 FC
83 27 C4 FD B3 07 F7 00 93 D7 17 40 23 2A F4 FC
83 27 44 FD 23 26 F4 FE 23 24 04 FE 6F 00 C0 0D
83 27 84 FD 23 22 F4 FE 23 20 04 FE 6F 00 40 0A
83 25 C4 FE 03 25 44 FE EF F0 1F E7 93 07 05 00
A3 09 F4 FC 83 27 80 4D 03 47 34 FD B7 06 00 01
93 86 F6 FF 33 77 D7 00 93 75 F7 0F 83 C6 D7 00
93 F6 06 00 13 86 06 00 93 86 05 00 B3 66 D6 00
A3 86 D7 00 93 56 87 00 93 F5 F6 0F 83 C6 E7 00
93 F6 06 00 13 86 06 00 93 86 05 00 B3 66 D6 00
23 87 D7 00 13 57 07 01 13 76 F7 0F 03 C7 F7 00
13 77 07 00 93 06 07 00 13 07 06 00 33 E7 E6 00
A3 87 E7 00 03 27 44 FE 83 27 C4 FD B3 07 F7 00
23 22 F4 FE 83 27 04 FE 93 87 17 00 23 20 F4 FE
03 27 04 FE 93 07 F0 27 E3 FC E7 F4 03 27 C4 FE
83 27 C4 FD B3 07 F7 00 23 26 F4 FE 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE 93 07 F0 1D
E3 F0 E7 F2 13 00 00 00 13 00 00 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 13 01 01 FE
23 2E 81 00 13 04 01 02 83 27 80 4D A3 89 07 00
23 26 04 FE 6F 00 00 0B 13 07 F0 0F 83 27 C4 FE
B3 07 F7 40 13 97 07 01 93 06 F0 0F 83 27 C4 FE
B3 87 F6 40 93 97 87 00 33 67 F7 00 93 06 F0 0F
83 27 C4 FE B3 87 F6 40 B3 66 F7 00 83 27 80 4D
37 07 00 01 13 07 F7 FF 33 F7 E6 00 93 75 F7 0F
83 C6 57 01 93 F6 06 00 13 86 06 00 93 86 05 00
B3 66 D6 00 A3 8A D7 00 93 56 87 00 93 F5 F6 0F
83 C6 67 01 93 F6 06 00 13 86 06 00 93 86 05 00
B3 66 D6 00 23 8B D7 00 13 57 07 01 13 76 F7 0F
03 C7 77 01 13 77 07 00 93 06 07 00 13 07 06 00
33 E7 E6 00 A3 8B E7 00 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE 93 07 E0 0F E3 F6 E7 F4
13 00 00 00 13 00 00 00 03 24 C1 01 13 01 01 02
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 83 27 80 4D 03 C7 37 00 13 67 07 F8
A3 81 E7 00 EF F0 9F EF 83 27 80 4D 03 C7 67 00
13 77 F7 01 23 83 E7 00 03 C7 77 00 13 77 07 00
A3 83 E7 00 83 27 80 4D 03 C7 A7 00 13 77 F7 03
23 85 E7 00 03 C7 B7 00 13 77 07 00 A3 85 E7 00
B7 07 00 FA 23 26 F4 FE B7 07 00 03 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 40 93 07 07 00
93 97 17 00 B3 87 E7 00 93 D7 27 40 23 22 F4 FE
83 27 44 FE 93 D7 17 40 B3 07 F0 40 23 20 F4 FE
83 27 44 FE 93 D7 17 40 23 2E F4 FC 83 26 C4 FD
03 26 04 FE 83 25 84 FE 03 25 C4 FE EF F0 DF CE
6F 00 00 00
@0000012B
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
34 FB FF FF 18 00 00 00 00 00 00 00
@00000136
00 00 00 80
