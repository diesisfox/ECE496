@00000000
00002197 A1418193 00010117 FF810113
00010433 0040006F
@00000006
000017B7 2147A683 FF010113 00112623
00100793 00F6A023 000017B7 DE878793
0006A823 40078613 0007A703 00478793
00E6AA23 FEC79AE3 4B8000EF 0000006F
02B507B3 02B51533 01A7D793 00651513
00F56533 00008067 80C1C683 01200793
04F68C63 000017B7 00269713 99C78793
00E787B3 0007A603 00001837 00001537
21C82303 21852883 00261713 00461793
00C70733 40C787B3 00571713 00379793
00670733 011787B3 00168693 20E82E23
20F52C23 80D18623 00008067 80C1C783
0C078A63 FFF78793 0FF7F793 80F18623
0C078463 00001737 99C70713 00279793
00F707B3 0007A683 000018B7 00001837
21882503 21C8A583 00269713 00469793
00D70733 40F68633 00571313 00361613
00771713 406585B3 00A60633 40D70733
02FC6537 20B8AE23 20C82C23 00B70733
66650513 00E55A63 D8100593 02B685B3
00A585B3 20B8AE23 40D787B3 00579793
40D787B3 035C6737 00C787B3 66670713
00F75A63 E2100793 02F686B3 00E68633
20C82C23 FA03A7B7 99A78793 00F5D463
20F8AE23 FCA3A7B7 99A78793 00F65463
20F82C23 00008067 FA03A7B7 00001737
99A78793 20F72E23 FCA3A7B7 00001737
99A78793 20F72C23 00008067 80C1C783
000015B7 2185A803 00279713 000017B7
99C78793 00E787B3 00257713 0007A783
0C070463 00679713 00E80833 2105AC23
000018B7 00157713 21C8A683 08070A63
00679713 00E686B3 20D8AE23 00279713
00F70733 00771713 40F70733 02FC6637
00D70733 66660613 00E65A63 D8100693
02D786B3 00C686B3 20D8AE23 00479713
40F70733 00571713 40F70733 035C6637
01070733 66660613 00E65A63 E2100713
02E787B3 00C78833 2105AC23 FA03A737
99A70713 00E6D463 20E8AE23 FCA3A737
99A70713 00E85463 20E5AC23 00008067
00857513 F6050CE3 00679713 40E686B3
20D8AE23 F69FF06F 00457713 F40702E3
00679713 40E80833 2105AC23 F35FF06F
00050E13 00000313 00000713 00000613
00000F93 00000813 00000793 00000693
10000E93 10000F37 02FF8FB3 00130313
41070733 01031313 01C70733 01035313
02C686B3 02C7B533 01F686B3 41F75F93
02C787B3 00A686B3 00669693 00070613
01A7D793 00F6E7B3 00179793 00B787B3
05D30063 02C60533 41F7D693 02C61733
01A55513 02F788B3 00671713 00A76733
02F79833 01A8D893 00681813 01186833
00E80533 F8AF52E3 0FF37513 00008067
00000513 00008067 80C1C783 FF010113
00812623 00279713 000017B7 99C78793
00E787B3 0007AF83 000017B7 2187A303
000017B7 21C7A403 000017B7 2147A283
00912423 1E000393 10000E13 10000EB7
00040893 28000F13 00000513 00000593
00000793 00000693 00000713 00000613
00000813 02F80833 40B70733 00150513
01051513 01170733 01055513 02C686B3
02C7B5B3 010686B3 41F75813 02C787B3
00B686B3 00669693 00070613 01A7D793
00F6E7B3 00179793 006787B3 07C50263
02C605B3 41F7D693 02C61733 01A5D593
00671713 00B76733 02F784B3 02F795B3
01A4D493 00659593 0095E5B3 00B704B3
F89ED2E3 00A2A623 FFFF0F13 01F888B3
F40F1CE3 FFF38393 01F30333 F40392E3
00C12403 00812483 01010113 00008067
00000513 00A2A623 FFFF0F13 01F888B3
F20F14E3 FD1FF06F 00100793 00D796B3
02D05E63 000017B7 2147A703 00000813
00B807B3 00F72423 00A72223 00000793
00178793 00C72623 0FF7F793 FED7CAE3
00180813 0FF87813 FCD84CE3 00008067
80C1C783 FD010113 01812623 00279713
000017B7 99C78793 00E787B3 0007A503
000017B7 2187A703 000017B7 21C7AC03
000017B7 2147A783 02812623 02912423
03212223 03312023 01412E23 01512C23
01612A23 01712823 01912423 01A12223
01B12023 00551F13 00070813 02000E93
10000893 10000337 28000F93 20000393
FE0E8293 000C0593 00000E13 00000413
00000613 00000693 00000A13 00000913
00000493 00000993 02D989B3 40C90633
00B60633 00140413 01041413 01045413
029A0A33 02D4B933 014989B3 02D486B3
00060493 01298633 00661613 41F4D993
01A6D693 00D666B3 00169693 010686B3
2F140A63 02948B33 41F6DA13 02949633
01AB5B13 00661613 01666933 02D68AB3
02D69633 01AADA93 00661613 01566633
00C90AB3 F95352E3 00028613 00C7A423
01C7A223 02000693 FFF68693 0087A623
0FF6F693 FE069AE3 00160613 FECE90E3
020E0E13 01E585B3 F3FE1AE3 020E8E93
01E80833 F07E9EE3 00400A13 10000393
10000437 1E000693 4146DAB3 28000693
4146D9B3 00100693 014512B3 014698B3
00070E13 00000913 01491EB3 00197493
000C0B13 00000B93 00C0006F 000F0B93
000F8B13 009BE6B3 001B8F13 01628FB3
FE0686E3 00000593 00000613 00000693
00000C93 00000D13 00000813 00000313
030C8CB3 40CD0633 01660633 00158593
01059593 0105D593 02D30333 0306BD33
006C8333 030686B3 00060813 01A30633
00661613 41F85313 01A6D693 00D666B3
00169693 01C686B3 1C758263 03080633
41F6DC93 03081D33 01A65613 006D1D13
00CD6D33 02D68DB3 02D69633 01ADDD93
00661613 01B66633 00CD0DB3 F9B452E3
014B9BB3 00000613 01D606B3 00D7A423
0177A223 00000693 00168693 00B7A623
0FF6F693 FF16CAE3 00160613 0FF67613
FD164CE3 F13F6CE3 00190913 005E0E33
EF591CE3 FFFA0A13 EC0A16E3 00000493
00100393 10000E13 10000EB7 28000413
1E000913 00000F13 0014F293 000C0313
005F66B3 0097A423 00650FB3 001F0F13
00069E63 0077A223 000F8313 005F66B3
00650FB3 001F0F13 FE0686E3 00000613
00000993 00000893 00000693 00000A93
00000813 00000A13 02DA0A33 40C98633
00660633 00188893 01089893 0108D893
030A8AB3 02D835B3 015A0A33 02D806B3
00060813 00BA0633 00661613 41F85A13
01A6D693 00D666B3 00169693 00E686B3
09C88A63 030805B3 41F6DA93 030819B3
01A5D593 00699993 00B9E9B3 02D68633
02D695B3 01A65613 00659593 00C5E633
00C985B3 F8BED2E3 0117A623 F48F16E3
00148493 00A70733 F1249EE3 02C12403
02812483 02412903 02012983 01C12A03
01812A83 01412B03 01012B83 00C12C03
00812C83 00412D03 00012D83 03010113
00008067 00000413 D41FF06F 00000593
E71FF06F 00000893 0117A623 EE8F16E3
FA1FF06F 000017B7 2147A603 FFF00593
0FF00793 00062823 01079713 00879693
00D76733 00F76733 00E62A23 FFF78793
FEB794E3 00008067 000017B7 2147A603
000016B7 99C68693 04C68793 00062823
44C68693 0007A703 00478793 00E62A23
FED79AE3 00008067 000017B7 2147A683
000017B7 DE878793 0006A823 40078613
0007A703 00478793 00E6AA23 FEC79AE3
00008067
@00000267
0003999A 0001CCCD 0000E666 00007333
0000399A 00001CCD 00000E66 00000733
0000039A 000001CD 000000E6 00000073
0000003A 0000001D 0000000E 00000007
00000004 00000002 00000001 009D4200
009D4300 009E4401 009E4401 009F4502
009F4602 00A04702 00A04803 00A14803
00A14904 00A14A04 00A24B04 00A24C05
00A34C05 00A34D05 00A44E06 00A44F06
00A44F07 00A55007 00A55107 00A65208
00A65308 00A75309 00A75409 00A85509
00A8560A 00A8570A 00A9570B 00A9580B
00AA590B 00AA5A0C 00AB5B0C 00AB5B0D
00AB5C0D 00AC5D0D 00AC5E0E 00AD5F0E
00AD5F0E 00AE600F 00AE610F 00AF6210
00AF6310 00AF6310 00B06411 00B06511
00B16612 00B16612 00B26712 00B26813
00B26913 00B36A14 00B36A14 00B46B14
00B46C15 00B56D15 00B56E16 00B66E16
00B66F16 00B67017 00B77117 00B77217
00B87218 00B87318 00B97419 00B97519
00BA7619 00BA761A 00BA771A 00BB781B
00BB791B 00BC791B 00BC7A1C 00BD7B1C
00BD7C1D 00BD7D1D 00BE7D1D 00BE7E1E
00BF7F1E 00BF801F 00C0811F 00C0811F
00C18220 00C18320 00C18420 00C28521
00C28621 00C38622 00C38722 00C48822
00C48923 00C58A23 00C58A24 00C58B24
00C68C24 00C68D25 00C78E25 00C78E26
00C88F26 00C89026 00C99127 00C99227
00C99228 00CA9328 00CA9428 00CB9529
00CB9629 00CC962A 00CC972A 00CD982A
00CD992B 00CD9A2B 00CE9A2C 00CE9B2C
00CF9C2C 00CF9D2D 00D09E2D 00D09F2E
00D19F2E 00D1A02E 00D2A12F 00D2A22F
00D2A330 00D3A330 00D3A430 00D4A531
00D4A631 00D5A732 00D5A732 00D6A832
00D6A933 00D7AA33 00D7AB34 00D7AC34
00D8AC34 00D8AD35 00D9AE35 00D9AF36
00DAB036 00DAB137 00DBB137 00DBB237
00DCB338 00DCB438 00DCB539 00DDB639
00DDB639 00DEB73A 00DEB83A 00DFB93B
00DFBA3B 00E0BA3B 00E0BB3C 00E1BC3C
00E1BD3D 00E1BE3D 00E2BF3D 00E2BF3E
00E3C03E 00E3C13F 00E4C23F 00E4C340
00E5C440 00E5C440 00E6C541 00E6C641
00E7C742 00E7C842 00E7C942 00E8C943
00E8CA43 00E9CB44 00E9CC44 00EACD44
00EACE45 00EBCF45 00EBCF46 00ECD046
00ECD147 00EDD247 00EDD347 00EED448
00EED448 00EED549 00EFD649 00EFD749
00F0D84A 00F0D94A 00F1D94B 00F1DA4B
00F2DB4C 00F2DC4C 00F3DD4C 00F3DE4D
00F4DF4D 00F4DF4E 00F5E04E 00F5E14E
00F5E24F 00F6E34F 00F6E450 00F7E550
00F7E551 00F8E651 00F8E751 00F9E852
00F9E952 00FAEA53 00FAEB53 00FBEB54
00FBEC54 00FCED54 00FCEE55 00FDEF55
00FDF056 00FEF056 00FEF156 00FEF257
00FFF357 00FFF45C 00FFF462 00FFF468
00FFF56D 00FFF572 00FFF677 00FFF67C
00FFF680 00FFF785 00FFF789 00FFF88E
00FFF892 00FFF896 00FFF99B 00FFF99F
00FFF9A2 00FFFAA7 00FFFAAA 00FFFAAE
00FFFAB2 00FFFBB6 00FFFBB9 00FFFBBD
00FFFCC1 00FFFCC4 00FFFCC7 00FFFCCB
00FFFDCE 00FFFDD2 00FFFDD5 00FFFDD8
00FFFEDB 00FFFEDE 00FFFEE2 00FFFFE5
00FFFFE8 00FFFFEB 00000000 00598DFC
005A8EFC 005B8FFC 005B90FC 005C91FC
005D91FC 005E92FC 005F93FC 005F94FC
006095FC 006196FC 006297FC 006398FC
006399FC 00649AFC 00659AFC 00669BFC
00679CFC 00679DFC 00689EFC 00699FFC
006AA0FC 006BA1FD 006BA2FD 006CA2FD
006DA3FD 006EA4FD 006FA5FD 006FA6FD
0070A7FD 0071A8FD 0072A9FD 0073AAFD
0073ABFD 0074ABFD 0075ACFD 0076ADFD
0077AEFD 0077AFFD 0078B0FD 0079B1FD
007AB2FD 007BB3FD 007BB3FD 007CB4FD
007DB5FD 007EB6FD 007FB7FD 007FB8FD
0080B9FD 0081BAFD 0082BBFD 0083BBFD
0083BCFD 0084BDFD 0085BEFD 0086BFFD
0087C0FD 0087C1FD 0088C2FD 0089C3FD
008AC4FD 008BC4FD 008BC5FD 008CC6FE
008DC7FE 008EC8FE 008FC9FE 008FCAFE
0090CBFE 0091CCFE 0092CCFE 0093CDFE
0093CEFE 0094CFFE 0095D0FE 0096D1FE
0097D2FE 0097D3FE 0098D4FE 0099D5FE
009AD5FE 009BD6FE 009BD7FE 009CD8FE
009DD9FE 009EDAFE 009FDBFE 009FDCFE
00A0DDFE 00A1DDFE 00A2DEFE 00A3DFFE
00A3E0FE 00A4E1FE 00A5E2FE 00A6E3FE
00A7E4FE 00A7E5FE 00A8E6FE 00A9E6FE
00AAE7FE 00ABE8FE 00ABE9FE 00ACEAFE
00ADEBFE 00AEECFE 00AFEDFF 00AFEEFF
00B0EEFF 00B1EFFF 00B2F0FF 00B3F1FF
00B3F2FF 00B4F3FF 00B5F4FF 00B6F5FF
00B7F6FF 00B7F7FF 00B8F7FF 00B9F8FF
00BAF9FF 00BBFAFF 00BBFBFF 00BCFCFF
00BDFDFF 00BEFEFF 00BFFFFF 00BFFFFF
00BEFFFE 00BEFEFD 00BEFEFC 00BDFEFB
00BDFDFB 00BDFDFA 00BCFDF9 00BCFCF8
00BCFCF7 00BBFCF7 00BBFBF6 00BBFBF5
00BAFBF4 00BAFAF3 00BAFAF3 00B9FAF2
00B9F9F1 00B9F9F0 00B8F9EF 00B8F8EF
00B8F8EE 00B7F8ED 00B7F7EC 00B7F7EB
00B6F7EB 00B6F6EA 00B6F6E9 00B5F6E8
00B5F5E7 00B5F5E7 00B4F5E6 00B4F4E5
00B4F4E4 00B3F4E3 00B3F3E3 00B3F3E2
00B2F3E1 00B2F2E0 00B2F2DF 00B1F2DF
00B1F1DE 00B1F1DD 00B0F1DC 00B0F0DB
00B0F0DB 00AFF0DA 00AFEFD9 00AFEFD8
00AEEFD7 00AEEED7 00AEEED6 00ADEED5
00ADEDD4 00ADEDD3 00ACEDD3 00ACECD2
00ACECD1 00ABECD0 00ABEBCF 00ABEBCF
00AAEBCE 00AAEACD 00AAEACC 00A9EACB
00A9E9CB 00A9E9CA 00A8E9C9 00A8E8C8
00A8E8C7 00A7E8C7 00A7E7C6 00A7E7C5
00A6E7C4 00A6E6C3 00A6E6C3 00A5E6C2
00A5E5C1 00A5E5C0 00A4E5BF 00A4E4BF
00A4E4BE 00A3E4BD 00A3E3BC 00A3E3BB
00A2E3BB 00A2E3BA 00A1E2B9 00A1E2B8
00A1E2B7 00A0E1B7 00A0E1B6 00A0E1B5
009FE0B4 009FE0B3 009FE0B3 009EDFB2
009EDFB1 009EDFB0 009DDEAF 009DDEAF
009DDEAE 009CDDAD 009CDDAC 009CDDAB
009BDCAB 009BDCAA 009BDCA9 009ADBA8
009ADBA7 009ADBA7 0099DAA6 0099DAA5
0099DAA4 0098D9A3 0098D9A3 0098D9A2
0097D8A1 0097D8A0 0097D89F 0096D79F
0096D79E 0096D79D 0095D69C 0095D69B
0095D69B 0094D59A 0094D599
@0000047A
00000014 00000000 00527A03 01017C01
07020D1B 00000001 00000010 0000001C
FFFFEDF8 00000018 00000000
@00000485
80000000 FCA3999A FA03999A
