@00000000
97 11 00 00 93 81 01 B8 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 40 00
@00000006
03 27 00 38 13 01 01 FF 23 26 11 00 83 47 37 00
37 05 00 01 93 06 F0 0F 93 E7 07 F8 A3 01 F7 00
13 05 F5 FF A3 09 07 00 13 96 06 01 93 97 86 00
B3 E7 C7 00 B3 E7 D7 00 B3 F7 A7 00 93 F5 F7 0F
13 D6 87 00 03 48 57 01 13 76 F6 0F A3 0A B7 00
83 45 67 01 93 D7 07 01 23 0B C7 00 03 46 77 01
93 F7 F7 0F A3 0B F7 00 93 86 F6 FF E3 9E 06 FA
83 47 67 00 B7 06 60 03 37 06 A0 FC 93 F7 F7 01
23 03 F7 00 83 47 77 00 A3 03 07 00 83 47 A7 00
B7 05 00 03 37 05 00 FA 93 F7 F7 03 23 05 F7 00
83 47 B7 00 A3 05 07 00 EF 00 80 0D 6F 00 00 00
B3 07 B5 02 33 15 B5 02 93 D7 A7 01 13 15 65 00
33 65 F5 00 67 80 00 00 13 0E 05 00 13 03 00 00
13 07 00 00 13 06 00 00 93 0F 00 00 13 08 00 00
93 07 00 00 93 06 00 00 93 0E 00 10 37 0F 00 10
B3 8F FF 02 13 03 13 00 33 07 07 41 13 13 03 01
33 07 C7 01 13 53 03 01 B3 86 C6 02 33 B5 C7 02
B3 86 F6 01 93 5F F7 41 B3 87 C7 02 B3 86 A6 00
93 96 66 00 13 06 07 00 93 D7 A7 01 B3 E7 F6 00
93 97 17 00 B3 87 B7 00 63 00 D3 05 33 05 C6 02
93 D6 F7 41 33 17 C6 02 13 55 A5 01 B3 88 F7 02
13 17 67 00 33 67 A7 00 33 98 F7 02 93 D8 A8 01
13 18 68 00 33 68 18 01 33 05 E8 00 E3 52 AF F8
13 75 F3 0F 67 80 00 00 13 05 00 00 67 80 00 00
B7 A2 01 00 B3 87 A5 40 93 82 A2 99 33 87 57 02
03 2F 00 38 13 01 01 FF B7 03 00 01 23 26 81 00
23 24 91 00 23 22 21 01 93 04 00 1E 13 0E 00 10
B3 92 57 02 13 57 A7 01 B7 0E 00 10 93 83 F3 FF
93 92 62 00 B3 E2 E2 00 13 D3 12 40 33 04 A3 00
33 03 C3 00 93 08 04 00 93 0F 00 28 13 05 00 00
93 05 00 00 93 07 00 00 93 06 00 00 13 07 00 00
13 06 00 00 13 08 00 00 33 08 F8 02 33 07 B7 40
13 05 15 00 13 15 05 01 33 07 17 01 13 55 05 01
B3 86 C6 02 B3 B5 C7 02 B3 86 06 01 13 58 F7 41
B3 87 C7 02 B3 86 B6 00 93 96 66 00 13 06 07 00
93 D7 A7 01 B3 E7 F6 00 93 97 17 00 B3 87 67 00
63 0A C5 09 B3 05 C6 02 93 D6 F7 41 33 17 C6 02
93 D5 A5 01 13 17 67 00 33 67 B7 00 33 89 F7 02
B3 95 F7 02 13 59 A9 01 93 95 65 00 B3 E5 25 01
33 09 B7 00 E3 D2 2E F9 33 75 75 00 13 77 F5 0F
93 57 85 00 83 46 DF 00 93 F7 F7 0F A3 06 EF 00
03 47 EF 00 13 55 05 01 23 07 FF 00 83 47 FF 00
13 75 F5 0F A3 07 AF 00 93 8F FF FF B3 88 58 00
E3 96 0F F2 93 84 F4 FF 33 03 53 00 E3 9C 04 F0
03 24 C1 00 83 24 81 00 03 29 41 00 13 01 01 01
67 80 00 00 13 05 00 00 6F F0 5F FA 03 27 00 38
37 05 00 01 93 06 F0 0F A3 09 07 00 13 05 F5 FF
13 96 06 01 93 97 86 00 B3 E7 C7 00 B3 E7 D7 00
B3 F7 A7 00 93 F5 F7 0F 13 D6 87 00 03 48 57 01
13 76 F6 0F A3 0A B7 00 83 45 67 01 93 D7 07 01
23 0B C7 00 03 46 77 01 93 F7 F7 0F A3 0B F7 00
93 86 F6 FF E3 9E 06 FA 67 80 00 00
@000000D5
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
8C FC FF FF 18 00 00 00 00 00 00 00
@000000E0
00 00 00 80
