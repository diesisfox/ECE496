@00000000
97 11 00 00 93 81 01 B6 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 40 00
@00000006
03 27 00 36 13 01 01 FF 23 26 11 00 83 47 37 00
37 05 00 01 93 06 F0 0F 93 E7 07 F8 A3 01 F7 00
13 05 F5 FF A3 09 07 00 13 96 06 01 93 97 86 00
B3 E7 C7 00 B3 E7 D7 00 B3 F7 A7 00 93 F5 F7 0F
13 D6 87 00 03 48 57 01 13 76 F6 0F A3 0A B7 00
83 45 67 01 93 D7 07 01 23 0B C7 00 03 46 77 01
93 F7 F7 0F A3 0B F7 00 93 86 F6 FF E3 9E 06 FA
83 47 67 00 B7 06 60 03 37 06 A0 FC 93 F7 F7 01
23 03 F7 00 83 47 77 00 A3 03 07 00 83 47 A7 00
B7 05 00 03 37 05 00 FA 93 F7 F7 03 23 05 F7 00
83 47 B7 00 A3 05 07 00 EF 00 C0 0B 6F 00 00 00
13 0E 05 00 13 08 00 00 13 07 00 00 93 08 00 00
13 06 00 00 13 03 00 00 13 05 00 00 B7 0E 00 10
13 0F F0 0F 6F 00 80 00 63 04 E5 09 93 56 57 00
13 17 B7 01 93 96 66 00 93 57 A7 01 B3 E7 F6 00
93 D6 F7 41 33 03 F3 02 33 08 18 41 33 07 C8 01
13 05 15 00 13 75 F5 0F B3 86 C6 02 33 B8 C7 02
B3 86 66 00 B3 87 C7 02 B3 86 06 01 93 96 66 00
93 D7 A7 01 B3 E7 F6 00 33 86 F5 00 B3 06 E7 02
13 53 F6 41 33 18 E7 02 93 D6 A6 01 B3 07 C6 02
13 18 68 00 33 68 D8 00 B3 18 C6 02 93 D7 A7 01
93 98 68 00 B3 E8 F8 00 B3 87 08 01 E3 DE FE F6
67 80 00 00 B7 A2 01 00 B3 87 A5 40 93 82 A2 99
B3 86 57 02 03 2F 00 36 13 01 01 FF B7 03 00 01
23 26 81 00 23 24 91 00 23 22 21 01 93 04 00 1E
37 0E 00 10 B3 92 57 02 93 D6 A6 01 93 0E F0 0F
93 83 F3 FF 93 92 62 00 B3 E2 D2 00 33 07 55 00
33 03 56 00 13 54 17 40 13 53 13 40 93 08 04 00
93 0F 00 28 13 08 00 00 93 05 00 00 13 09 00 00
13 07 00 00 13 05 00 00 13 06 00 00 6F 00 80 00
63 0A D8 0D 93 56 57 00 13 17 B7 01 93 96 66 00
93 57 A7 01 B3 E7 F6 00 93 D6 F7 41 33 09 F9 02
33 06 A6 40 33 07 16 01 13 08 18 00 13 78 F8 0F
B3 86 B6 02 33 B6 B7 02 B3 86 26 01 B3 87 B7 02
B3 86 C6 00 93 96 66 00 93 D7 A7 01 B3 E7 F6 00
B3 05 F3 00 B3 06 E7 02 13 D9 F5 41 33 16 E7 02
93 D6 A6 01 B3 87 B5 02 13 16 66 00 33 66 D6 00
33 95 B5 02 93 D7 A7 01 13 15 65 00 33 65 F5 00
B3 07 A6 00 E3 5E FE F6 33 78 78 00 13 78 F8 0F
83 47 DF 00 A3 06 0F 01 83 47 EF 00 23 07 0F 00
83 47 FF 00 93 8F FF FF A3 07 0F 00 B3 88 58 00
E3 9A 0F F2 93 84 F4 FF 33 03 53 00 E3 90 04 F2
03 24 C1 00 83 24 81 00 03 29 41 00 13 01 01 01
67 80 00 00 13 08 F0 0F 6F F0 5F FB 03 27 00 36
37 05 00 01 93 06 F0 0F A3 09 07 00 13 05 F5 FF
13 96 06 01 93 97 86 00 B3 E7 C7 00 B3 E7 D7 00
B3 F7 A7 00 93 F5 F7 0F 13 D6 87 00 03 48 57 01
13 76 F6 0F A3 0A B7 00 83 45 67 01 93 D7 07 01
23 0B C7 00 03 46 77 01 93 F7 F7 0F A3 0B F7 00
93 86 F6 FF E3 9E 06 FA 67 80 00 00
@000000CD
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
AC FC FF FF 18 00 00 00 00 00 00 00
@000000D8
00 00 00 80
