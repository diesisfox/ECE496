@00000000
97 21 00 00 93 81 41 A1 17 01 01 00 13 01 81 FF
33 04 01 00 6F 00 40 00
@00000018
B7 17 00 00 83 A6 47 21 13 01 01 FF 23 26 11 00
93 07 10 00 23 A0 F6 00 B7 17 00 00 93 87 87 DE
23 A8 06 00 13 86 07 40 03 A7 07 00 93 87 47 00
23 AA E6 00 E3 9A C7 FE EF 00 80 4B 6F 00 00 00
B3 07 B5 02 33 15 B5 02 93 D7 A7 01 13 15 65 00
33 65 F5 00 67 80 00 00 83 C6 C1 80 93 07 20 01
63 8C F6 04 B7 17 00 00 13 97 26 00 93 87 C7 99
B3 87 E7 00 03 A6 07 00 37 18 00 00 37 15 00 00
03 23 C8 21 83 28 85 21 13 17 26 00 93 17 46 00
33 07 C7 00 B3 87 C7 40 13 17 57 00 93 97 37 00
33 07 67 00 B3 87 17 01 93 86 16 00 23 2E E8 20
23 2C F5 20 23 86 D1 80 67 80 00 00 83 C7 C1 80
63 8A 07 0C 93 87 F7 FF 93 F7 F7 0F 23 86 F1 80
63 84 07 0C 37 17 00 00 13 07 C7 99 93 97 27 00
B3 07 F7 00 83 A6 07 00 B7 18 00 00 37 18 00 00
03 25 88 21 83 A5 C8 21 13 97 26 00 93 97 46 00
33 07 D7 00 33 86 F6 40 13 13 57 00 13 16 36 00
13 17 77 00 B3 85 65 40 33 06 A6 00 33 07 D7 40
37 65 FC 02 23 AE B8 20 23 2C C8 20 33 07 B7 00
13 05 65 66 63 5A E5 00 93 05 10 D8 B3 85 B6 02
B3 85 A5 00 23 AE B8 20 B3 87 D7 40 93 97 57 00
B3 87 D7 40 37 67 5C 03 B3 87 C7 00 13 07 67 66
63 5A F7 00 93 07 10 E2 B3 86 F6 02 33 86 E6 00
23 2C C8 20 B7 A7 03 FA 93 87 A7 99 63 D4 F5 00
23 AE F8 20 B7 A7 A3 FC 93 87 A7 99 63 54 F6 00
23 2C F8 20 67 80 00 00 B7 A7 03 FA 37 17 00 00
93 87 A7 99 23 2E F7 20 B7 A7 A3 FC 37 17 00 00
93 87 A7 99 23 2C F7 20 67 80 00 00 83 C7 C1 80
B7 15 00 00 03 A8 85 21 13 97 27 00 B7 17 00 00
93 87 C7 99 B3 87 E7 00 13 77 25 00 83 A7 07 00
63 04 07 0C 13 97 67 00 33 08 E8 00 23 AC 05 21
B7 18 00 00 13 77 15 00 83 A6 C8 21 63 0A 07 08
13 97 67 00 B3 86 E6 00 23 AE D8 20 13 97 27 00
33 07 F7 00 13 17 77 00 33 07 F7 40 37 66 FC 02
33 07 D7 00 13 06 66 66 63 5A E6 00 93 06 10 D8
B3 86 D7 02 B3 86 C6 00 23 AE D8 20 13 97 47 00
33 07 F7 40 13 17 57 00 33 07 F7 40 37 66 5C 03
33 07 07 01 13 06 66 66 63 5A E6 00 13 07 10 E2
B3 87 E7 02 33 88 C7 00 23 AC 05 21 37 A7 03 FA
13 07 A7 99 63 D4 E6 00 23 AE E8 20 37 A7 A3 FC
13 07 A7 99 63 54 E8 00 23 AC E5 20 67 80 00 00
13 75 85 00 E3 0C 05 F6 13 97 67 00 B3 86 E6 40
23 AE D8 20 6F F0 9F F6 13 77 45 00 E3 02 07 F4
13 97 67 00 33 08 E8 40 23 AC 05 21 6F F0 5F F3
13 0E 05 00 13 03 00 00 13 07 00 00 13 06 00 00
93 0F 00 00 13 08 00 00 93 07 00 00 93 06 00 00
93 0E 00 10 37 0F 00 10 B3 8F FF 02 13 03 13 00
33 07 07 41 13 13 03 01 33 07 C7 01 13 53 03 01
B3 86 C6 02 33 B5 C7 02 B3 86 F6 01 93 5F F7 41
B3 87 C7 02 B3 86 A6 00 93 96 66 00 13 06 07 00
93 D7 A7 01 B3 E7 F6 00 93 97 17 00 B3 87 B7 00
63 00 D3 05 33 05 C6 02 93 D6 F7 41 33 17 C6 02
13 55 A5 01 B3 88 F7 02 13 17 67 00 33 67 A7 00
33 98 F7 02 93 D8 A8 01 13 18 68 00 33 68 18 01
33 05 E8 00 E3 52 AF F8 13 75 F3 0F 67 80 00 00
13 05 00 00 67 80 00 00 83 C7 C1 80 13 01 01 FF
23 26 81 00 13 97 27 00 B7 17 00 00 93 87 C7 99
B3 87 E7 00 83 AF 07 00 B7 17 00 00 03 A3 87 21
B7 17 00 00 03 A4 C7 21 B7 17 00 00 83 A2 47 21
23 24 91 00 93 03 00 1E 13 0E 00 10 B7 0E 00 10
93 08 04 00 13 0F 00 28 13 05 00 00 93 05 00 00
93 07 00 00 93 06 00 00 13 07 00 00 13 06 00 00
13 08 00 00 33 08 F8 02 33 07 B7 40 13 05 15 00
13 15 05 01 33 07 17 01 13 55 05 01 B3 86 C6 02
B3 B5 C7 02 B3 86 06 01 13 58 F7 41 B3 87 C7 02
B3 86 B6 00 93 96 66 00 13 06 07 00 93 D7 A7 01
B3 E7 F6 00 93 97 17 00 B3 87 67 00 63 02 C5 07
B3 05 C6 02 93 D6 F7 41 33 17 C6 02 93 D5 A5 01
13 17 67 00 33 67 B7 00 B3 84 F7 02 B3 95 F7 02
93 D4 A4 01 93 95 65 00 B3 E5 95 00 B3 04 B7 00
E3 D2 9E F8 23 A6 A2 00 13 0F FF FF B3 88 F8 01
E3 1C 0F F4 93 83 F3 FF 33 03 F3 01 E3 92 03 F4
03 24 C1 00 83 24 81 00 13 01 01 01 67 80 00 00
13 05 00 00 23 A6 A2 00 13 0F FF FF B3 88 F8 01
E3 14 0F F2 6F F0 1F FD 93 07 10 00 B3 96 D7 00
63 5E D0 02 B7 17 00 00 03 A7 47 21 13 08 00 00
B3 07 B8 00 23 24 F7 00 23 22 A7 00 93 07 00 00
93 87 17 00 23 26 C7 00 93 F7 F7 0F E3 CA D7 FE
13 08 18 00 13 78 F8 0F E3 4C D8 FC 67 80 00 00
83 C7 C1 80 13 01 01 FD 23 26 81 01 13 97 27 00
B7 17 00 00 93 87 C7 99 B3 87 E7 00 03 A5 07 00
B7 17 00 00 03 A7 87 21 B7 17 00 00 03 AC C7 21
B7 17 00 00 83 A7 47 21 23 26 81 02 23 24 91 02
23 22 21 03 23 20 31 03 23 2E 41 01 23 2C 51 01
23 2A 61 01 23 28 71 01 23 24 91 01 23 22 A1 01
23 20 B1 01 13 1F 55 00 13 08 07 00 93 0E 00 02
93 08 00 10 37 03 00 10 93 0F 00 28 93 03 00 20
93 82 0E FE 93 05 0C 00 13 0E 00 00 13 04 00 00
13 06 00 00 93 06 00 00 13 0A 00 00 13 09 00 00
93 04 00 00 93 09 00 00 B3 89 D9 02 33 06 C9 40
33 06 B6 00 13 04 14 00 13 14 04 01 13 54 04 01
33 0A 9A 02 33 B9 D4 02 B3 89 49 01 B3 86 D4 02
93 04 06 00 33 86 29 01 13 16 66 00 93 D9 F4 41
93 D6 A6 01 B3 66 D6 00 93 96 16 00 B3 86 06 01
63 0A 14 2F 33 8B 94 02 13 DA F6 41 33 96 94 02
13 5B AB 01 13 16 66 00 33 69 66 01 B3 8A D6 02
33 96 D6 02 93 DA AA 01 13 16 66 00 33 66 56 01
B3 0A C9 00 E3 52 53 F9 13 86 02 00 23 A4 C7 00
23 A2 C7 01 93 06 00 02 93 86 F6 FF 23 A6 87 00
93 F6 F6 0F E3 9A 06 FE 13 06 16 00 E3 90 CE FE
13 0E 0E 02 B3 85 E5 01 E3 1A FE F3 93 8E 0E 02
33 08 E8 01 E3 9E 7E F0 13 0A 40 00 93 03 00 10
37 04 00 10 93 06 00 1E B3 DA 46 41 93 06 00 28
B3 D9 46 41 93 06 10 00 B3 12 45 01 B3 98 46 01
13 0E 07 00 13 09 00 00 B3 1E 49 01 93 74 19 00
13 0B 0C 00 93 0B 00 00 6F 00 C0 00 93 0B 0F 00
13 8B 0F 00 B3 E6 9B 00 13 8F 1B 00 B3 8F 62 01
E3 86 06 FE 93 05 00 00 13 06 00 00 93 06 00 00
93 0C 00 00 13 0D 00 00 13 08 00 00 13 03 00 00
B3 8C 0C 03 33 06 CD 40 33 06 66 01 93 85 15 00
93 95 05 01 93 D5 05 01 33 03 D3 02 33 BD 06 03
33 83 6C 00 B3 86 06 03 13 08 06 00 33 06 A3 01
13 16 66 00 13 53 F8 41 93 D6 A6 01 B3 66 D6 00
93 96 16 00 B3 86 C6 01 63 82 75 1C 33 06 08 03
93 DC F6 41 33 1D 08 03 13 56 A6 01 13 1D 6D 00
33 6D CD 00 B3 8D D6 02 33 96 D6 02 93 DD AD 01
13 16 66 00 33 66 B6 01 B3 0D CD 00 E3 52 B4 F9
B3 9B 4B 01 13 06 00 00 B3 06 D6 01 23 A4 D7 00
23 A2 77 01 93 06 00 00 93 86 16 00 23 A6 B7 00
93 F6 F6 0F E3 CA 16 FF 13 06 16 00 13 76 F6 0F
E3 4C 16 FD E3 6C 3F F1 13 09 19 00 33 0E 5E 00
E3 1C 59 EF 13 0A FA FF E3 16 0A EC 93 04 00 00
93 03 10 00 13 0E 00 10 B7 0E 00 10 13 04 00 28
13 09 00 1E 13 0F 00 00 93 F2 14 00 13 03 0C 00
B3 66 5F 00 23 A4 97 00 B3 0F 65 00 13 0F 1F 00
63 9E 06 00 23 A2 77 00 13 83 0F 00 B3 66 5F 00
B3 0F 65 00 13 0F 1F 00 E3 86 06 FE 13 06 00 00
93 09 00 00 93 08 00 00 93 06 00 00 93 0A 00 00
13 08 00 00 13 0A 00 00 33 0A DA 02 33 86 C9 40
33 06 66 00 93 88 18 00 93 98 08 01 93 D8 08 01
B3 8A 0A 03 B3 35 D8 02 33 0A 5A 01 B3 06 D8 02
13 08 06 00 33 06 BA 00 13 16 66 00 13 5A F8 41
93 D6 A6 01 B3 66 D6 00 93 96 16 00 B3 86 E6 00
63 8A C8 09 B3 05 08 03 93 DA F6 41 B3 19 08 03
93 D5 A5 01 93 99 69 00 B3 E9 B9 00 33 86 D6 02
B3 95 D6 02 13 56 A6 01 93 95 65 00 33 E6 C5 00
B3 85 C9 00 E3 D2 BE F8 23 A6 17 01 E3 16 8F F4
93 84 14 00 33 07 A7 00 E3 9E 24 F1 03 24 C1 02
83 24 81 02 03 29 41 02 83 29 01 02 03 2A C1 01
83 2A 81 01 03 2B 41 01 83 2B 01 01 03 2C C1 00
83 2C 81 00 03 2D 41 00 83 2D 01 00 13 01 01 03
67 80 00 00 13 04 00 00 6F F0 1F D4 93 05 00 00
6F F0 1F E7 93 08 00 00 23 A6 17 01 E3 16 8F EE
6F F0 1F FA B7 17 00 00 03 A6 47 21 93 05 F0 FF
93 07 F0 0F 23 28 06 00 13 97 07 01 93 96 87 00
33 67 D7 00 33 67 F7 00 23 2A E6 00 93 87 F7 FF
E3 94 B7 FE 67 80 00 00 B7 17 00 00 03 A6 47 21
B7 16 00 00 93 86 C6 99 93 87 C6 04 23 28 06 00
93 86 C6 44 03 A7 07 00 93 87 47 00 23 2A E6 00
E3 9A D7 FE 67 80 00 00 B7 17 00 00 83 A6 47 21
B7 17 00 00 93 87 87 DE 23 A8 06 00 13 86 07 40
03 A7 07 00 93 87 47 00 23 AA E6 00 E3 9A C7 FE
67 80 00 00
@0000099C
9A 99 03 00 CD CC 01 00 66 E6 00 00 33 73 00 00
9A 39 00 00 CD 1C 00 00 66 0E 00 00 33 07 00 00
9A 03 00 00 CD 01 00 00 E6 00 00 00 73 00 00 00
3A 00 00 00 1D 00 00 00 0E 00 00 00 07 00 00 00
04 00 00 00 02 00 00 00 01 00 00 00 00 42 9D 00
00 43 9D 00 01 44 9E 00 01 44 9E 00 02 45 9F 00
02 46 9F 00 02 47 A0 00 03 48 A0 00 03 48 A1 00
04 49 A1 00 04 4A A1 00 04 4B A2 00 05 4C A2 00
05 4C A3 00 05 4D A3 00 06 4E A4 00 06 4F A4 00
07 4F A4 00 07 50 A5 00 07 51 A5 00 08 52 A6 00
08 53 A6 00 09 53 A7 00 09 54 A7 00 09 55 A8 00
0A 56 A8 00 0A 57 A8 00 0B 57 A9 00 0B 58 A9 00
0B 59 AA 00 0C 5A AA 00 0C 5B AB 00 0D 5B AB 00
0D 5C AB 00 0D 5D AC 00 0E 5E AC 00 0E 5F AD 00
0E 5F AD 00 0F 60 AE 00 0F 61 AE 00 10 62 AF 00
10 63 AF 00 10 63 AF 00 11 64 B0 00 11 65 B0 00
12 66 B1 00 12 66 B1 00 12 67 B2 00 13 68 B2 00
13 69 B2 00 14 6A B3 00 14 6A B3 00 14 6B B4 00
15 6C B4 00 15 6D B5 00 16 6E B5 00 16 6E B6 00
16 6F B6 00 17 70 B6 00 17 71 B7 00 17 72 B7 00
18 72 B8 00 18 73 B8 00 19 74 B9 00 19 75 B9 00
19 76 BA 00 1A 76 BA 00 1A 77 BA 00 1B 78 BB 00
1B 79 BB 00 1B 79 BC 00 1C 7A BC 00 1C 7B BD 00
1D 7C BD 00 1D 7D BD 00 1D 7D BE 00 1E 7E BE 00
1E 7F BF 00 1F 80 BF 00 1F 81 C0 00 1F 81 C0 00
20 82 C1 00 20 83 C1 00 20 84 C1 00 21 85 C2 00
21 86 C2 00 22 86 C3 00 22 87 C3 00 22 88 C4 00
23 89 C4 00 23 8A C5 00 24 8A C5 00 24 8B C5 00
24 8C C6 00 25 8D C6 00 25 8E C7 00 26 8E C7 00
26 8F C8 00 26 90 C8 00 27 91 C9 00 27 92 C9 00
28 92 C9 00 28 93 CA 00 28 94 CA 00 29 95 CB 00
29 96 CB 00 2A 96 CC 00 2A 97 CC 00 2A 98 CD 00
2B 99 CD 00 2B 9A CD 00 2C 9A CE 00 2C 9B CE 00
2C 9C CF 00 2D 9D CF 00 2D 9E D0 00 2E 9F D0 00
2E 9F D1 00 2E A0 D1 00 2F A1 D2 00 2F A2 D2 00
30 A3 D2 00 30 A3 D3 00 30 A4 D3 00 31 A5 D4 00
31 A6 D4 00 32 A7 D5 00 32 A7 D5 00 32 A8 D6 00
33 A9 D6 00 33 AA D7 00 34 AB D7 00 34 AC D7 00
34 AC D8 00 35 AD D8 00 35 AE D9 00 36 AF D9 00
36 B0 DA 00 37 B1 DA 00 37 B1 DB 00 37 B2 DB 00
38 B3 DC 00 38 B4 DC 00 39 B5 DC 00 39 B6 DD 00
39 B6 DD 00 3A B7 DE 00 3A B8 DE 00 3B B9 DF 00
3B BA DF 00 3B BA E0 00 3C BB E0 00 3C BC E1 00
3D BD E1 00 3D BE E1 00 3D BF E2 00 3E BF E2 00
3E C0 E3 00 3F C1 E3 00 3F C2 E4 00 40 C3 E4 00
40 C4 E5 00 40 C4 E5 00 41 C5 E6 00 41 C6 E6 00
42 C7 E7 00 42 C8 E7 00 42 C9 E7 00 43 C9 E8 00
43 CA E8 00 44 CB E9 00 44 CC E9 00 44 CD EA 00
45 CE EA 00 45 CF EB 00 46 CF EB 00 46 D0 EC 00
47 D1 EC 00 47 D2 ED 00 47 D3 ED 00 48 D4 EE 00
48 D4 EE 00 49 D5 EE 00 49 D6 EF 00 49 D7 EF 00
4A D8 F0 00 4A D9 F0 00 4B D9 F1 00 4B DA F1 00
4C DB F2 00 4C DC F2 00 4C DD F3 00 4D DE F3 00
4D DF F4 00 4E DF F4 00 4E E0 F5 00 4E E1 F5 00
4F E2 F5 00 4F E3 F6 00 50 E4 F6 00 50 E5 F7 00
51 E5 F7 00 51 E6 F8 00 51 E7 F8 00 52 E8 F9 00
52 E9 F9 00 53 EA FA 00 53 EB FA 00 54 EB FB 00
54 EC FB 00 54 ED FC 00 55 EE FC 00 55 EF FD 00
56 F0 FD 00 56 F0 FE 00 56 F1 FE 00 57 F2 FE 00
57 F3 FF 00 5C F4 FF 00 62 F4 FF 00 68 F4 FF 00
6D F5 FF 00 72 F5 FF 00 77 F6 FF 00 7C F6 FF 00
80 F6 FF 00 85 F7 FF 00 89 F7 FF 00 8E F8 FF 00
92 F8 FF 00 96 F8 FF 00 9B F9 FF 00 9F F9 FF 00
A2 F9 FF 00 A7 FA FF 00 AA FA FF 00 AE FA FF 00
B2 FA FF 00 B6 FB FF 00 B9 FB FF 00 BD FB FF 00
C1 FC FF 00 C4 FC FF 00 C7 FC FF 00 CB FC FF 00
CE FD FF 00 D2 FD FF 00 D5 FD FF 00 D8 FD FF 00
DB FE FF 00 DE FE FF 00 E2 FE FF 00 E5 FF FF 00
E8 FF FF 00 EB FF FF 00 00 00 00 00 FC 8D 59 00
FC 8E 5A 00 FC 8F 5B 00 FC 90 5B 00 FC 91 5C 00
FC 91 5D 00 FC 92 5E 00 FC 93 5F 00 FC 94 5F 00
FC 95 60 00 FC 96 61 00 FC 97 62 00 FC 98 63 00
FC 99 63 00 FC 9A 64 00 FC 9A 65 00 FC 9B 66 00
FC 9C 67 00 FC 9D 67 00 FC 9E 68 00 FC 9F 69 00
FC A0 6A 00 FD A1 6B 00 FD A2 6B 00 FD A2 6C 00
FD A3 6D 00 FD A4 6E 00 FD A5 6F 00 FD A6 6F 00
FD A7 70 00 FD A8 71 00 FD A9 72 00 FD AA 73 00
FD AB 73 00 FD AB 74 00 FD AC 75 00 FD AD 76 00
FD AE 77 00 FD AF 77 00 FD B0 78 00 FD B1 79 00
FD B2 7A 00 FD B3 7B 00 FD B3 7B 00 FD B4 7C 00
FD B5 7D 00 FD B6 7E 00 FD B7 7F 00 FD B8 7F 00
FD B9 80 00 FD BA 81 00 FD BB 82 00 FD BB 83 00
FD BC 83 00 FD BD 84 00 FD BE 85 00 FD BF 86 00
FD C0 87 00 FD C1 87 00 FD C2 88 00 FD C3 89 00
FD C4 8A 00 FD C4 8B 00 FD C5 8B 00 FE C6 8C 00
FE C7 8D 00 FE C8 8E 00 FE C9 8F 00 FE CA 8F 00
FE CB 90 00 FE CC 91 00 FE CC 92 00 FE CD 93 00
FE CE 93 00 FE CF 94 00 FE D0 95 00 FE D1 96 00
FE D2 97 00 FE D3 97 00 FE D4 98 00 FE D5 99 00
FE D5 9A 00 FE D6 9B 00 FE D7 9B 00 FE D8 9C 00
FE D9 9D 00 FE DA 9E 00 FE DB 9F 00 FE DC 9F 00
FE DD A0 00 FE DD A1 00 FE DE A2 00 FE DF A3 00
FE E0 A3 00 FE E1 A4 00 FE E2 A5 00 FE E3 A6 00
FE E4 A7 00 FE E5 A7 00 FE E6 A8 00 FE E6 A9 00
FE E7 AA 00 FE E8 AB 00 FE E9 AB 00 FE EA AC 00
FE EB AD 00 FE EC AE 00 FF ED AF 00 FF EE AF 00
FF EE B0 00 FF EF B1 00 FF F0 B2 00 FF F1 B3 00
FF F2 B3 00 FF F3 B4 00 FF F4 B5 00 FF F5 B6 00
FF F6 B7 00 FF F7 B7 00 FF F7 B8 00 FF F8 B9 00
FF F9 BA 00 FF FA BB 00 FF FB BB 00 FF FC BC 00
FF FD BD 00 FF FE BE 00 FF FF BF 00 FF FF BF 00
FE FF BE 00 FD FE BE 00 FC FE BE 00 FB FE BD 00
FB FD BD 00 FA FD BD 00 F9 FD BC 00 F8 FC BC 00
F7 FC BC 00 F7 FC BB 00 F6 FB BB 00 F5 FB BB 00
F4 FB BA 00 F3 FA BA 00 F3 FA BA 00 F2 FA B9 00
F1 F9 B9 00 F0 F9 B9 00 EF F9 B8 00 EF F8 B8 00
EE F8 B8 00 ED F8 B7 00 EC F7 B7 00 EB F7 B7 00
EB F7 B6 00 EA F6 B6 00 E9 F6 B6 00 E8 F6 B5 00
E7 F5 B5 00 E7 F5 B5 00 E6 F5 B4 00 E5 F4 B4 00
E4 F4 B4 00 E3 F4 B3 00 E3 F3 B3 00 E2 F3 B3 00
E1 F3 B2 00 E0 F2 B2 00 DF F2 B2 00 DF F2 B1 00
DE F1 B1 00 DD F1 B1 00 DC F1 B0 00 DB F0 B0 00
DB F0 B0 00 DA F0 AF 00 D9 EF AF 00 D8 EF AF 00
D7 EF AE 00 D7 EE AE 00 D6 EE AE 00 D5 EE AD 00
D4 ED AD 00 D3 ED AD 00 D3 ED AC 00 D2 EC AC 00
D1 EC AC 00 D0 EC AB 00 CF EB AB 00 CF EB AB 00
CE EB AA 00 CD EA AA 00 CC EA AA 00 CB EA A9 00
CB E9 A9 00 CA E9 A9 00 C9 E9 A8 00 C8 E8 A8 00
C7 E8 A8 00 C7 E8 A7 00 C6 E7 A7 00 C5 E7 A7 00
C4 E7 A6 00 C3 E6 A6 00 C3 E6 A6 00 C2 E6 A5 00
C1 E5 A5 00 C0 E5 A5 00 BF E5 A4 00 BF E4 A4 00
BE E4 A4 00 BD E4 A3 00 BC E3 A3 00 BB E3 A3 00
BB E3 A2 00 BA E3 A2 00 B9 E2 A1 00 B8 E2 A1 00
B7 E2 A1 00 B7 E1 A0 00 B6 E1 A0 00 B5 E1 A0 00
B4 E0 9F 00 B3 E0 9F 00 B3 E0 9F 00 B2 DF 9E 00
B1 DF 9E 00 B0 DF 9E 00 AF DE 9D 00 AF DE 9D 00
AE DE 9D 00 AD DD 9C 00 AC DD 9C 00 AB DD 9C 00
AB DC 9B 00 AA DC 9B 00 A9 DC 9B 00 A8 DB 9A 00
A7 DB 9A 00 A7 DB 9A 00 A6 DA 99 00 A5 DA 99 00
A4 DA 99 00 A3 D9 98 00 A3 D9 98 00 A2 D9 98 00
A1 D8 97 00 A0 D8 97 00 9F D8 97 00 9F D7 96 00
9E D7 96 00 9D D7 96 00 9C D6 95 00 9B D6 95 00
9B D6 95 00 9A D5 94 00 99 D5 94 00
@000011E8
14 00 00 00 00 00 00 00 03 7A 52 00 01 7C 01 01
1B 0D 02 07 01 00 00 00 10 00 00 00 1C 00 00 00
F8 ED FF FF 18 00 00 00 00 00 00 00
@00001214
00 00 00 80 9A 99 A3 FC 9A 99 03 FA
