@00000000
00001197 07C18193 00010117 FF810113
00010433 7AC0006F
@00000006
FE010113 00812E23 02010413 FEA42623
FEB42423 FEC42583 00058813 41F5D593
00058893 FE842583 00058613 41F5D593
00058693 02C88533 030685B3 00B505B3
02C80533 02C837B3 00050713 00F586B3
00068793 00679693 01A75313 0066E333
41A7D393 00030793 00078513 01C12403
02010113 00008067 FE010113 00812E23
02010413 80C1C703 01200793 08F70863
80C1C783 00078693 000017B7 80478713
00269793 00F707B3 0007A783 FEF42623
FEC42703 00070793 00279793 00E787B3
00579793 00078713 000017B7 87C7A783
00F70733 000017B7 86E7AE23 FEC42703
00070793 00479793 40E787B3 00379793
00078713 000017B7 8807A783 00F70733
000017B7 88E7A023 80C1C783 00178793
0FF7F713 80E18623 0080006F 00000013
01C12403 02010113 00008067 FE010113
00812E23 02010413 80C1C783 1A078263
80C1C783 FFF78793 0FF7F713 80E18623
80C1C783 02079463 000017B7 FA03A737
99A70713 86E7AE23 000017B7 FCA3A737
99A70713 88E7A023 16C0006F 80C1C783
00078693 000017B7 80478713 00269793
00F707B3 0007A783 FEF42623 FEC42703
00070793 00279793 00E787B3 00579793
40F00733 000017B7 87C7A783 00F70733
000017B7 86E7AE23 FEC42703 00070793
00471713 40E787B3 00379793 00078713
000017B7 8807A783 00F70733 000017B7
88E7A023 FEC42703 00070793 00279793
00E787B3 00779793 40E78733 000017B7
87C7A783 00F70733 02FC67B7 66678793
02E7D263 FEC42703 D8100793 02F70733
02FC67B7 66678793 00F70733 000017B7
86E7AE23 FEC42703 00070793 00479793
40E787B3 00579793 40E78733 000017B7
8807A783 00F70733 035C67B7 66678793
02E7D263 FEC42703 E2100793 02F70733
035C67B7 66678793 00F70733 000017B7
88E7A023 000017B7 87C7A703 FA03A7B7
99A78793 00F75A63 000017B7 FA03A737
99A70713 86E7AE23 000017B7 8807A703
FCA3A7B7 99A78793 00F75E63 000017B7
FCA3A737 99A70713 88E7A023 0080006F
00000013 01C12403 02010113 00008067
FD010113 02812623 03010413 00050793
FCF40FA3 80C1C783 00078693 000017B7
80478713 00269793 00F707B3 0007A783
FEF42623 FDF44783 0027F793 02078263
FEC42783 00679713 000017B7 8807A783
00F70733 000017B7 88E7A023 02C0006F
FDF44783 0047F793 02078063 000017B7
8807A703 FEC42783 00679793 40F70733
000017B7 88E7A023 FDF44783 0017F793
02078263 FEC42783 00679713 000017B7
87C7A783 00F70733 000017B7 86E7AE23
02C0006F FDF44783 0087F793 02078063
000017B7 87C7A703 FEC42783 00679793
40F70733 000017B7 86E7AE23 FEC42703
00070793 00279793 00E787B3 00779793
40E78733 000017B7 87C7A783 00F70733
02FC67B7 66678793 02E7D263 FEC42703
D8100793 02F70733 02FC67B7 66678793
00F70733 000017B7 86E7AE23 FEC42703
00070793 00479793 40E787B3 00579793
40E78733 000017B7 8807A783 00F70733
035C67B7 66678793 02E7D263 FEC42703
E2100793 02F70733 035C67B7 66678793
00F70733 000017B7 88E7A023 000017B7
87C7A703 FA03A7B7 99A78793 00F75A63
000017B7 FA03A737 99A70713 86E7AE23
000017B7 8807A703 FCA3A7B7 99A78793
00F75A63 000017B7 FCA3A737 99A70713
88E7A023 00000013 02C12403 03010113
00008067 FC010113 02112E23 02812C23
04010413 FCA42623 FCB42423 0FF00793
FEF41223 FE042623 FE042423 FE041323
08C0006F FEC42583 FEC42503 B05FF0EF
FEA42023 FE842583 FE842503 AF5FF0EF
FCA42E23 FE042703 FDC42783 00F70733
100007B7 06E7C463 FE042703 FDC42783
40F707B3 FCC42703 00F707B3 FCF42C23
FE842583 FEC42503 AB9FF0EF 00050793
00179793 FC842703 00F707B3 FCF42A23
FD842783 FEF42623 FD442783 FEF42423
FE645783 00178793 FEF41323 FE645703
FE445783 F6E7F8E3 0080006F 00000013
FE645783 0FF7F793 00078513 03C12083
03812403 04010113 00008067 FD010113
02112623 02812423 03010413 80C1C783
00078693 000017B7 80478713 00269793
00F707B3 0007A783 FCF42E23 000017B7
8807A783 FEF42623 FE042423 0800006F
000017B7 87C7A783 FEF42223 FE042023
0440006F FEC42583 FE442503 EB9FF0EF
00050793 FCF40DA3 000017B7 8847A783
FDB44703 00E7A623 FE442703 FDC42783
00F707B3 FEF42223 FE042783 00178793
FEF42023 FE042703 27F00793 FAE7FCE3
FEC42703 FDC42783 00F707B3 FEF42623
FE842783 00178793 FEF42423 FE842703
1DF00793 F6E7FEE3 00000013 00000013
02C12083 02812403 03010113 00008067
FE010113 00812E23 02010413 000017B7
8847A783 0007A823 FE042623 0500006F
0FF00713 FEC42783 40F707B3 01079713
0FF00693 FEC42783 40F687B3 00879793
00F766B3 0FF00713 FEC42783 40F70733
000017B7 8847A783 00E6E733 00E7AA23
FEC42783 00178793 FEF42623 FEC42703
0FE00793 FAE7F6E3 00000013 00000013
01C12403 02010113 00008067 FE010113
00812E23 02010413 000017B7 8847A783
0007A823 FE042623 0500006F 0FF00713
FEC42783 40F707B3 01079713 0FF00693
FEC42783 40F687B3 00879793 00F766B3
0FF00713 FEC42783 40F70733 000017B7
8847A783 00E6E733 00E7AA23 FEC42783
00178793 FEF42623 FEC42703 0FE00793
FAE7F6E3 00000013 00000013 01C12403
02010113 00008067 FF010113 00112623
00812423 01010413 000017B7 8847A783
00100713 00E7A023 EC9FF0EF 000017B7
8847A783 0007A223 000017B7 8847A783
0007A423 DC9FF0EF 0000006F
@00000201
0003999A 0001CCCD 0000E666 00007333
0000399A 00001CCD 00000E66 00000733
0000039A 000001CD 000000E6 00000073
0000003A 0000001D 0000000E 00000007
00000004 00000002 00000001
@00000214
00000014 00000000 00527A03 01017C01
07020D1B 00000001 00000010 0000001C
FFFFF790 00000018 00000000
@0000021F
FA03999A FCA3999A 80000000
