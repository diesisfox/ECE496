`include "../AXI5-Lite.sv"

module ip_gpio_main (
    ports
);
    
endmodule
