@00000000
00003197 48818193 00010117 FF810113
00010433 0040006F
@00000006
000037B7 C8C7A603 FF010113 000017B7
BF078793 00112623 00100713 06C78593
00E62023 46878793 0007A683 00078713
FFC78793 00D62A23 FEE598E3 6BC000EF
FE051EE3 50C000EF FE051AE3 504000EF
FE050AE3 FE9FF06F 02B507B3 02B51533
01A7D793 00651513 00F56533 00008067
8141C683 01200793 04F68A63 000017B7
00269713 BF078793 00E787B3 0007A603
00003537 80C1A303 C9052883 00261713
00461793 00C70733 40C787B3 00571713
00379793 00670733 011787B3 00168693
80E1A623 C8F52823 80D18A23 00008067
8141C783 0C078863 FFF78793 0FF7F793
80F18A23 0C078263 00001737 BF070713
00279793 00F707B3 0007A683 00003837
C9082503 80C1A583 00269713 00469793
00D70733 40F68633 00571313 00361613
00771713 406585B3 00A60633 40D70733
02FC6537 80B1A623 C8C82823 00B70733
66650513 00E55A63 D8100593 02B685B3
00A585B3 80B1A623 40D787B3 00579793
40D787B3 035C6737 00C787B3 66670713
00F75A63 E2100793 02F686B3 00E68633
C8C82823 FA03A7B7 99A78793 00F5D463
80F1A623 FCA3A7B7 99A78793 00F65463
C8F82823 00008067 FA03A7B7 99A78793
80F1A623 FCA3A7B7 00003737 99A78793
C8F72823 00008067 8141C783 000035B7
C905A803 00279713 000017B7 BF078793
00E787B3 00257713 0007A783 0C070263
00679713 00E80833 C905A823 00157713
80C1A683 08070A63 00679713 00E686B3
80D1A623 00279713 00F70733 00771713
40F70733 02FC6637 00D70733 66660613
00E65A63 D8100693 02D786B3 00C686B3
80D1A623 00479713 40F70733 00571713
40F70733 035C6637 01070733 66660613
00E65A63 E2100713 02E787B3 00C78833
C905A823 FA03A737 99A70713 00E6D463
80E1A623 FCA3A737 99A70713 00E85463
C8E5A823 00008067 00857513 F6050CE3
00679713 40E686B3 80D1A623 F69FF06F
00457713 F40704E3 00679713 40E80833
C905A823 F39FF06F 00050E13 00000313
00000713 00000613 00000F93 00000813
00000793 00000693 0FF00E93 10000F37
02FF8FB3 00130313 41070733 01031313
01C70733 01035313 02C686B3 02C7B533
01F686B3 41F75F93 02C787B3 00A686B3
00669693 00070613 01A7D793 00F6E7B3
00179793 00B787B3 05D30063 02C60533
41F7D693 02C61733 01A55513 02F788B3
00671713 00A76733 02F79833 01A8D893
00681813 01186833 00E80533 F8AF52E3
0FF37513 00008067 0FF00513 00008067
8141C783 FF010113 00812623 00279713
000017B7 BF078793 00E787B3 0007AF83
000037B7 C907A303 80C1A403 000037B7
C8C7A283 00912423 1E000393 0FF00E13
10000EB7 00040893 28000F13 00000513
00000593 00000793 00000693 00000713
00000613 00000813 02F80833 40B70733
00150513 01051513 01170733 01055513
02C686B3 02C7B5B3 010686B3 41F75813
02C787B3 00B686B3 00669693 00070613
01A7D793 00F6E7B3 00179793 006787B3
07C50263 02C605B3 41F7D693 02C61733
01A5D593 00671713 00B76733 02F784B3
02F795B3 01A4D493 00659593 0095E5B3
00B704B3 F89ED2E3 00A2A623 FFFF0F13
01F888B3 F40F1CE3 FFF38393 01F30333
F40392E3 00C12403 00812483 01010113
00008067 0FF00513 00A2A623 FFFF0F13
01F888B3 F20F14E3 FD1FF06F 00100793
00D796B3 02D05E63 000037B7 C8C7A703
00000813 00B807B3 00F72423 00A72223
00000793 00178793 00C72623 0FF7F793
FED7CAE3 00180813 0FF87813 FCD84CE3
00008067 00155793 00279713 000017B7
BF078793 00E787B3 00157513 00003737
04C7A783 C8C72683 00050E63 40078613
0007A703 00478793 00E6AA23 FEF61AE3
00008067 3FC78713 00072583 00070613
FFC70713 00B6AA23 FEC798E3 00008067
000037B7 C887A703 FF010113 01212023
00912223 8101A783 00072483 00112623
00812423 00000513 08978C63 FFF7C793
0097F433 00F47793 0A079263 01047793
06078263 8141C683 01200793 00100513
04F68A63 000017B7 00269713 BF078793
00E787B3 0007A603 00003837 80C1AE03
C9082303 00261713 00461793 00C70733
40C787B3 00571713 00379793 01C70733
006787B3 00168693 80E1A623 C8F82823
80D18A23 02047413 0A041663 8101A783
00F4C7B3 0067D793 00F7F793 02079C63
00C12083 00812403 8091A823 00412483
00012903 01010113 00008067 00078513
B99FF0EF 01047793 00100513 FA078CE3
F55FF06F 0064D793 0FF7F793 00179693
01C6F713 000016B7 BF068693 00E686B3
0017F713 04C6A783 000036B7 C8C6A683
04070A63 40078613 0007A703 00478793
00E6AA23 FEF61AE3 00C12083 00812403
8091A823 00412483 00012903 01010113
00008067 A2DFF0EF 8101A783 00100513
00F4C7B3 0067D793 00F7F793 F4078AE3
F85FF06F 3FC78713 00072583 00070613
FFC70713 00B6AA23 FEC798E3 00C12083
00812403 8091A823 00412483 00012903
01010113 00008067 8141C783 FB010113
05212023 00279713 000017B7 BF078793
00E787B3 0007A783 00003737 C9072903
03412C23 03612823 03712623 03812423
04112623 04812423 04912223 03312E23
03512A23 03912223 03A12023 01B12E23
00F12023 00579C13 02000B13 00000513
10000A37 00003BB7 80C1A483 FE0B0D13
00000A93 0FF00993 00001CB7 00000413
00000613 00000793 00000813 00000713
00000693 00000593 02F585B3 40C70733
00970733 00140413 01041413 01045413
02D80833 02F6B633 010585B3 02F687B3
00070693 00C58733 00671713 41F6D593
01A7D793 00F767B3 00179793 012787B3
37340E63 02D68633 41F7D813 02D69733
01A65613 00671713 00C76733 02F788B3
02F79633 01A8D893 00661613 01166633
00C708B3 F91A52E3 00040793 00F50533
2EACC863 C8CBA783 000D0693 00D7A423
0157A223 02000713 FFF70713 0087A623
0FF77713 FE071AE3 00168693 FEDB10E3
020A8A93 28000713 018484B3 F2EA90E3
020B0B13 20000713 01890933 EEEB1EE3
00400C13 0FF00993 10000A37 00003737
C9072903 00012703 00000593 1E000893
01871CB3 28000813 000C0713 00100413
4188D8B3 41885833 01841433 001C9D13
00058C13 00070593 80C1A483 00080713
00BC1B33 001C7D93 000C0813 009C84B3
00100A93 00001337 00070C13 00C0006F
009D04B3 001A8A93 FFFA8E93 01DDE733
419484B3 FE0706E3 00000E13 00000693
00000713 00000F93 00000293 00000613
00000F13 02EF0F33 40D286B3 009686B3
001E0E13 010E1E13 010E5E13 02CF8FB3
02E632B3 01FF0F33 02E60733 00068613
005F06B3 00669693 41F65F13 01A75713
00E6E733 00171713 01270733 233E0A63
02C606B3 41F75F93 02C612B3 01A6D693
00629293 00D2E2B3 02E703B3 02E716B3
01A3D393 00669693 0076E6B3 00D283B3
F87A52E3 000E0693 00BE9EB3 00000613
01660733 00E7A423 01D7A223 00000713
00170713 00D7A623 0FF77713 FE874AE3
00160613 0FF67613 FC864CE3 01C50533
18A34A63 F18AE6E3 000C0713 00080C13
001C0C13 00070813 01990933 ED1C16E3
FFF58C13 E80C14E3 00012C83 00003737
C9072483 00000A93 00100D13 10000937
001C9B13 01812023 80C1A403 0157A423
001AFD93 01940433 00100A13 0FF00993
00001837 28000C13 0100006F 01A7A223
008B0433 001A0A13 FFFA0713 01B76733
41940433 FE0704E3 00000693 00000E93
00000593 00000713 00000E13 00000613
00000313 02E30333 40DE86B3 008686B3
00158593 01059593 0105D593 02CE0E33
02E63EB3 01C30333 02E60733 00068613
01D306B3 00669693 41F65313 01A75713
00E6E733 00171713 00970733 11358463
02C606B3 41F75E13 02C61EB3 01A6D693
006E9E93 00DEEEB3 02E70F33 02E716B3
01AF5F13 00669693 01E6E6B3 00DE8F33
F9E952E3 00058713 00B50533 00E7A623
08A84E63 0B8A0463 C8CBA783 F35FF06F
A41FF0EF D00508E3 00100C13 04C12083
04812403 04412483 04012903 03C12983
03812A03 03412A83 03012B03 02C12B83
02412C83 02012D03 01C12D83 000C0513
02812C03 05010113 00008067 0FF00793
CBDFF06F 00B12623 01112423 01012223
9E1FF0EF FA0512E3 C8CBA783 00C12583
00812883 00412803 00001337 E49FF06F
0FF00693 0FF00E13 E01FF06F 9B5FF0EF
00001837 F6051AE3 F78A10E3 001A8A93
1E000793 019484B3 00FA8C63 C8CBA783
E59FF06F 0FF00713 0FF00593 F2DFF06F
00012C03 F49FF06F
@000002FC
0003999A 0001CCCD 0000E666 00007333
0000399A 00001CCD 00000E66 00000733
0000039A 000001CD 000000E6 00000073
0000003A 0000001D 0000000E 00000007
00000004 00000002 00000001 0000105C
0000145C 0000185C 00001C5C 0000205C
0000245C 00000C5C 0000285C 00640700
00660901 00670A01 00690C02 006A0D02
006C0F03 006E1003 006F1204 00711404
00731505 00741705 00761806 00771A06
00791B07 007B1D07 007C1F08 007E2008
007F2209 00812309 0083250A 0084260A
0086280B 00882A0B 00892B0C 008B2D0C
008C2E0D 008E300D 0090310E 0091330E
0093340F 0094360F 00963810 00983910
00993B11 009B3C11 009D3E12 009E3F12
00A04113 00A14313 00A34414 00A54614
00A64715 00A84915 00A94A16 00AB4C16
00AD4E17 00AE4F17 00B05118 00B25218
00B35419 00B55519 00B6571A 00B8591A
00BA5A1B 00BB5C1B 00BD5D1C 00BE5F1C
00C0601D 00C2621D 00C3641E 00C5651E
00C7671F 00C8681F 00CA6A20 00CB6C21
00CC6E24 00CD7027 00CE732A 00CE752E
00CF7731 00D07A34 00D17C37 00D27E3B
00D3803E 00D38341 00D48544 00D58747
00D68A4B 00D78C4E 00D78E51 00D89154
00D99357 00DA955B 00DB985E 00DC9A61
00DC9C64 00DD9F68 00DEA16B 00DFA36E
00E0A671 00E0A874 00E1AA78 00E2AD7B
00E3AF7E 00E4B181 00E4B484 00E5B688
00E6B88B 00E7BB8E 00E8BD91 00E9BF95
00E9C198 00EAC49B 00EBC69E 00ECC8A1
00EDCBA5 00EDCDA8 00EECFAB 00EFD2AE
00F0D4B2 00F1D6B5 00F2D9B8 00F2DBBB
00F3DDBE 00F4E0C2 00F5E2C5 00F6E4C8
00F6E7CB 00F7E9CE 00F8EBD2 00F9EED5
00FAF0D8 00FBF2DB 00FBF5DF 00FCF7E2
00FDF9E5 00FEFCE8 00FFFEEB 00FDFEED
00F9FDED 00F5FCEE 00F1FAEE 00EDF9EE
00E9F8EF 00E5F6EF 00E1F5EF 00DDF4EF
00D9F2F0 00D5F1F0 00D1F0F0 00CDEEF1
00C9EDF1 00C5ECF1 00C1EAF1 00BDE9F2
00B9E8F2 00B5E6F2 00B1E5F3 00ADE4F3
00A9E2F3 00A5E1F3 00A1E0F4 009DDEF4
0099DDF4 0095DCF4 0091DAF5 008DD9F5
0089D8F5 0085D6F6 0081D5F6 007DD4F6
0079D2F6 0075D1F7 0071D0F7 006DCEF7
0069CDF8 0065CCF8 0061CAF8 005DC9F8
0059C8F9 0055C6F9 0051C5F9 004DC4FA
0049C2FA 0045C1FA 0041C0FA 003DBEFB
0039BDFB 0035BCFB 0031BAFC 002DB9FC
0029B8FC 0025B6FC 0021B5FD 001DB4FD
0019B2FD 0015B1FE 0011B0FE 000DAEFE
0009ADFE 0005ACFF 0001AAFF 0000A8FC
0000A5F8 0000A3F4 0000A0F0 00009DEC
00009BE8 000098E4 000096E0 000093DC
000090D8 00008ED4 00008BD0 000088CC
000086C8 000083C4 000080C0 00007EBC
00007BB8 000079B4 000076B0 000073AC
000071A8 00006EA4 00006BA0 0000699C
00006698 00006494 00006190 00005E8C
00005C88 00005984 00005680 0000547C
00005178 00004E74 00004C70 0000496C
00004768 00004464 00004160 00003F5C
00003C58 00003954 00003750 0000344C
00003148 00002F44 00002C40 00002A3C
00002738 00002434 00002230 00001F2C
00001C28 00001A24 00001720 0000141C
00001218 00000F14 00000D10 00000A0C
00000708 00000504 00000200 00FFFFFF
00FEFEFE 00FDFDFD 00FCFCFC 00FBFBFB
00FAFAFA 00F9F9F9 00F8F8F8 00F7F7F7
00F6F6F6 00F5F5F5 00F4F4F4 00F3F3F3
00F2F2F2 00F1F1F1 00F0F0F0 00EFEFEF
00EEEEEE 00EDEDED 00ECECEC 00EBEBEB
00EAEAEA 00E9E9E9 00E8E8E8 00E7E7E7
00E6E6E6 00E5E5E5 00E4E4E4 00E3E3E3
00E2E2E2 00E1E1E1 00E0E0E0 00DFDFDF
00DEDEDE 00DDDDDD 00DCDCDC 00DBDBDB
00DADADA 00D9D9D9 00D8D8D8 00D7D7D7
00D6D6D6 00D5D5D5 00D4D4D4 00D3D3D3
00D2D2D2 00D1D1D1 00D0D0D0 00CFCFCF
00CECECE 00CDCDCD 00CCCCCC 00CBCBCB
00CACACA 00C9C9C9 00C8C8C8 00C7C7C7
00C6C6C6 00C5C5C5 00C4C4C4 00C3C3C3
00C2C2C2 00C1C1C1 00C0C0C0 00BFBFBF
00BEBEBE 00BDBDBD 00BCBCBC 00BBBBBB
00BABABA 00B9B9B9 00B8B8B8 00B7B7B7
00B6B6B6 00B5B5B5 00B4B4B4 00B3B3B3
00B2B2B2 00B1B1B1 00B0B0B0 00AFAFAF
00AEAEAE 00ADADAD 00ACACAC 00ABABAB
00AAAAAA 00A9A9A9 00A8A8A8 00A7A7A7
00A6A6A6 00A5A5A5 00A4A4A4 00A3A3A3
00A2A2A2 00A1A1A1 00A0A0A0 009F9F9F
009E9E9E 009D9D9D 009C9C9C 009B9B9B
009A9A9A 00999999 00989898 00979797
00969696 00959595 00949494 00939393
00929292 00919191 00909090 008F8F8F
008E8E8E 008D8D8D 008C8C8C 008B8B8B
008A8A8A 00898989 00888888 00878787
00868686 00858585 00848484 00838383
00828282 00818181 00808080 007F7F7F
007E7E7E 007D7D7D 007C7C7C 007B7B7B
007A7A7A 00797979 00787878 00777777
00767676 00757575 00747474 00737373
00727272 00717171 00707070 006F6F6F
006E6E6E 006D6D6D 006C6C6C 006B6B6B
006A6A6A 00696969 00686868 00676767
00666666 00656565 00646464 00636363
00626262 00616161 00606060 005F5F5F
005E5E5E 005D5D5D 005C5C5C 005B5B5B
005A5A5A 00595959 00585858 00575757
00565656 00555555 00545454 00535353
00525252 00515151 00505050 004F4F4F
004E4E4E 004D4D4D 004C4C4C 004B4B4B
004A4A4A 00494949 00484848 00474747
00464646 00454545 00444444 00434343
00424242 00414141 00404040 003F3F3F
003E3E3E 003D3D3D 003C3C3C 003B3B3B
003A3A3A 00393939 00383838 00373737
00363636 00353535 00343434 00333333
00323232 00313131 00303030 002F2F2F
002E2E2E 002D2D2D 002C2C2C 002B2B2B
002A2A2A 00292929 00282828 00272727
00262626 00252525 00242424 00232323
00222222 00212121 00202020 001F1F1F
001E1E1E 001D1D1D 001C1C1C 001B1B1B
001A1A1A 00191919 00181818 00171717
00161616 00151515 00141414 00131313
00121212 00111111 00101010 000F0F0F
000E0E0E 000D0D0D 000C0C0C 000B0B0B
000A0A0A 00090909 00080808 00070707
00060606 00050505 00040404 00030303
00020202 00010101 00000000 009D4200
009D4300 009E4401 009E4401 009F4502
009F4602 00A04702 00A04803 00A14803
00A14904 00A14A04 00A24B04 00A24C05
00A34C05 00A34D05 00A44E06 00A44F06
00A44F07 00A55007 00A55107 00A65208
00A65308 00A75309 00A75409 00A85509
00A8560A 00A8570A 00A9570B 00A9580B
00AA590B 00AA5A0C 00AB5B0C 00AB5B0D
00AB5C0D 00AC5D0D 00AC5E0E 00AD5F0E
00AD5F0E 00AE600F 00AE610F 00AF6210
00AF6310 00AF6310 00B06411 00B06511
00B16612 00B16612 00B26712 00B26813
00B26913 00B36A14 00B36A14 00B46B14
00B46C15 00B56D15 00B56E16 00B66E16
00B66F16 00B67017 00B77117 00B77217
00B87218 00B87318 00B97419 00B97519
00BA7619 00BA761A 00BA771A 00BB781B
00BB791B 00BC791B 00BC7A1C 00BD7B1C
00BD7C1D 00BD7D1D 00BE7D1D 00BE7E1E
00BF7F1E 00BF801F 00C0811F 00C0811F
00C18220 00C18320 00C18420 00C28521
00C28621 00C38622 00C38722 00C48822
00C48923 00C58A23 00C58A24 00C58B24
00C68C24 00C68D25 00C78E25 00C78E26
00C88F26 00C89026 00C99127 00C99227
00C99228 00CA9328 00CA9428 00CB9529
00CB9629 00CC962A 00CC972A 00CD982A
00CD992B 00CD9A2B 00CE9A2C 00CE9B2C
00CF9C2C 00CF9D2D 00D09E2D 00D09F2E
00D19F2E 00D1A02E 00D2A12F 00D2A22F
00D2A330 00D3A330 00D3A430 00D4A531
00D4A631 00D5A732 00D5A732 00D6A832
00D6A933 00D7AA33 00D7AB34 00D7AC34
00D8AC34 00D8AD35 00D9AE35 00D9AF36
00DAB036 00DAB137 00DBB137 00DBB237
00DCB338 00DCB438 00DCB539 00DDB639
00DDB639 00DEB73A 00DEB83A 00DFB93B
00DFBA3B 00E0BA3B 00E0BB3C 00E1BC3C
00E1BD3D 00E1BE3D 00E2BF3D 00E2BF3E
00E3C03E 00E3C13F 00E4C23F 00E4C340
00E5C440 00E5C440 00E6C541 00E6C641
00E7C742 00E7C842 00E7C942 00E8C943
00E8CA43 00E9CB44 00E9CC44 00EACD44
00EACE45 00EBCF45 00EBCF46 00ECD046
00ECD147 00EDD247 00EDD347 00EED448
00EED448 00EED549 00EFD649 00EFD749
00F0D84A 00F0D94A 00F1D94B 00F1DA4B
00F2DB4C 00F2DC4C 00F3DD4C 00F3DE4D
00F4DF4D 00F4DF4E 00F5E04E 00F5E14E
00F5E24F 00F6E34F 00F6E450 00F7E550
00F7E551 00F8E651 00F8E751 00F9E852
00F9E952 00FAEA53 00FAEB53 00FBEB54
00FBEC54 00FCED54 00FCEE55 00FDEF55
00FDF056 00FEF056 00FEF156 00FEF257
00FFF357 00FFF45C 00FFF462 00FFF468
00FFF56D 00FFF572 00FFF677 00FFF67C
00FFF680 00FFF785 00FFF789 00FFF88E
00FFF892 00FFF896 00FFF99B 00FFF99F
00FFF9A2 00FFFAA7 00FFFAAA 00FFFAAE
00FFFAB2 00FFFBB6 00FFFBB9 00FFFBBD
00FFFCC1 00FFFCC4 00FFFCC7 00FFFCCB
00FFFDCE 00FFFDD2 00FFFDD5 00FFFDD8
00FFFEDB 00FFFEDE 00FFFEE2 00FFFFE5
00FFFFE8 00FFFFEB 00FFFFEE 00598DFC
005A8EFC 005B8FFC 005B90FC 005C91FC
005D91FC 005E92FC 005F93FC 005F94FC
006095FC 006196FC 006297FC 006398FC
006399FC 00649AFC 00659AFC 00669BFC
00679CFC 00679DFC 00689EFC 00699FFC
006AA0FC 006BA1FD 006BA2FD 006CA2FD
006DA3FD 006EA4FD 006FA5FD 006FA6FD
0070A7FD 0071A8FD 0072A9FD 0073AAFD
0073ABFD 0074ABFD 0075ACFD 0076ADFD
0077AEFD 0077AFFD 0078B0FD 0079B1FD
007AB2FD 007BB3FD 007BB3FD 007CB4FD
007DB5FD 007EB6FD 007FB7FD 007FB8FD
0080B9FD 0081BAFD 0082BBFD 0083BBFD
0083BCFD 0084BDFD 0085BEFD 0086BFFD
0087C0FD 0087C1FD 0088C2FD 0089C3FD
008AC4FD 008BC4FD 008BC5FD 008CC6FE
008DC7FE 008EC8FE 008FC9FE 008FCAFE
0090CBFE 0091CCFE 0092CCFE 0093CDFE
0093CEFE 0094CFFE 0095D0FE 0096D1FE
0097D2FE 0097D3FE 0098D4FE 0099D5FE
009AD5FE 009BD6FE 009BD7FE 009CD8FE
009DD9FE 009EDAFE 009FDBFE 009FDCFE
00A0DDFE 00A1DDFE 00A2DEFE 00A3DFFE
00A3E0FE 00A4E1FE 00A5E2FE 00A6E3FE
00A7E4FE 00A7E5FE 00A8E6FE 00A9E6FE
00AAE7FE 00ABE8FE 00ABE9FE 00ACEAFE
00ADEBFE 00AEECFE 00AFEDFF 00AFEEFF
00B0EEFF 00B1EFFF 00B2F0FF 00B3F1FF
00B3F2FF 00B4F3FF 00B5F4FF 00B6F5FF
00B7F6FF 00B7F7FF 00B8F7FF 00B9F8FF
00BAF9FF 00BBFAFF 00BBFBFF 00BCFCFF
00BDFDFF 00BEFEFF 00BFFFFF 00BFFFFF
00BEFFFE 00BEFEFD 00BEFEFC 00BDFEFB
00BDFDFB 00BDFDFA 00BCFDF9 00BCFCF8
00BCFCF7 00BBFCF7 00BBFBF6 00BBFBF5
00BAFBF4 00BAFAF3 00BAFAF3 00B9FAF2
00B9F9F1 00B9F9F0 00B8F9EF 00B8F8EF
00B8F8EE 00B7F8ED 00B7F7EC 00B7F7EB
00B6F7EB 00B6F6EA 00B6F6E9 00B5F6E8
00B5F5E7 00B5F5E7 00B4F5E6 00B4F4E5
00B4F4E4 00B3F4E3 00B3F3E3 00B3F3E2
00B2F3E1 00B2F2E0 00B2F2DF 00B1F2DF
00B1F1DE 00B1F1DD 00B0F1DC 00B0F0DB
00B0F0DB 00AFF0DA 00AFEFD9 00AFEFD8
00AEEFD7 00AEEED7 00AEEED6 00ADEED5
00ADEDD4 00ADEDD3 00ACEDD3 00ACECD2
00ACECD1 00ABECD0 00ABEBCF 00ABEBCF
00AAEBCE 00AAEACD 00AAEACC 00A9EACB
00A9E9CB 00A9E9CA 00A8E9C9 00A8E8C8
00A8E8C7 00A7E8C7 00A7E7C6 00A7E7C5
00A6E7C4 00A6E6C3 00A6E6C3 00A5E6C2
00A5E5C1 00A5E5C0 00A4E5BF 00A4E4BF
00A4E4BE 00A3E4BD 00A3E3BC 00A3E3BB
00A2E3BB 00A2E3BA 00A1E2B9 00A1E2B8
00A1E2B7 00A0E1B7 00A0E1B6 00A0E1B5
009FE0B4 009FE0B3 009FE0B3 009EDFB2
009EDFB1 009EDFB0 009DDEAF 009DDEAF
009DDEAE 009CDDAD 009CDDAC 009CDDAB
009BDCAB 009BDCAA 009BDCA9 009ADBA8
009ADBA7 009ADBA7 0099DAA6 0099DAA5
0099DAA4 0098D9A3 0098D9A3 0098D9A2
0097D8A1 0097D8A0 0097D89F 0096D79F
0096D79E 0096D79D 0095D69C 0095D69B
0095D69B 0094D59A 0094D599 00CCFFFF
00CCFEFE 00CBFEFC 00CBFDFB 00CAFDF9
00CAFCF8 00CAFCF6 00C9FBF5 00C9FAF3
00C9FAF2 00C8F9F0 00C8F9EF 00C7F8ED
00C7F7EC 00C7F7EA 00C6F6E9 00C6F6E7
00C6F5E6 00C5F5E4 00C5F4E3 00C4F3E2
00C4F3E0 00C4F2DF 00C3F2DD 00C3F1DC
00C3F0DA 00C2F0D9 00C2EFD7 00C1EFD6
00C1EED4 00C1EED3 00C0EDD1 00C0ECD0
00C0ECCE 00BFEBCD 00BFEBCB 00BEEACA
00BEEAC8 00BEE9C7 00BDE8C5 00BDE8C4
00BDE7C3 00BCE7C1 00BCE6C0 00BBE5BE
00BBE5BD 00BBE4BB 00BAE4BA 00BAE3B8
00BAE3B7 00B9E2B5 00B9E1B4 00B8E1B2
00B8E0B1 00B8E0AF 00B7DFAE 00B7DEAC
00B7DEAB 00B6DDA9 00B6DDA8 00B5DCA7
00B5DCA5 00B5DBA4 00B4DAA2 00B4DAA1
00B4D99F 00B5D99E 00B5D89C 00B5D89B
00B5D799 00B6D698 00B6D696 00B6D595
00B6D593 00B7D492 00B7D490 00B7D38F
00B7D38D 00B8D28C 00B8D18A 00B8D189
00B8D087 00B9D086 00B9CF84 00B9CF83
00B9CE81 00BACD7F 00BACD7E 00BACC7C
00BACC7B 00BBCB79 00BBCB78 00BBCA76
00BBC975 00BCC973 00BCC872 00BCC870
00BCC76F 00BDC76D 00BDC66C 00BDC66A
00BDC569 00BEC467 00BEC466 00BEC364
00BEC363 00BFC261 00BFC260 00BFC15E
00BFC05D 00C0C05B 00C0BF5A 00C0BF58
00C0BE57 00C1BE55 00C1BD54 00C1BC52
00C1BC51 00C2BB4F 00C2BB4E 00C2BA4C
00C2BA4B 00C3B949 00C3B948 00C3B846
00C3B745 00C4B743 00C4B642 00C4B641
00C4B541 00C4B440 00C3B340 00C3B240
00C3B13F 00C3B03F 00C3B03F 00C2AF3E
00C2AE3E 00C2AD3E 00C2AC3D 00C2AB3D
00C1AA3D 00C1A93C 00C1A93C 00C1A83C
00C1A73B 00C1A63B 00C0A53B 00C0A43A
00C0A33A 00C0A33A 00C0A239 00BFA139
00BFA039 00BF9F38 00BF9E38 00BF9D38
00BE9D37 00BE9C37 00BE9B37 00BE9A36
00BE9936 00BE9836 00BD9735 00BD9735
00BD9635 00BD9534 00BD9434 00BC9334
00BC9233 00BC9133 00BC9033 00BC9032
00BB8F32 00BB8E32 00BB8D31 00BB8C31
00BB8B31 00BA8A30 00BA8A30 00BA8930
00BA882F 00BA872F 00BA862F 00B9852E
00B9842E 00B9842E 00B9832D 00B9822D
00B8812D 00B8802C 00B87F2C 00B87E2C
00B77D2C 00B67C2C 00B67B2C 00B5792B
00B5782B 00B4772B 00B4762B 00B3752B
00B2742B 00B2722B 00B1712B 00B1702B
00B06F2A 00B06E2A 00AF6C2A 00AF6B2A
00AE6A2A 00AD692A 00AD682A 00AC672A
00AC652A 00AB642A 00AB6329 00AA6229
00A96129 00A96029 00A85E29 00A85D29
00A75C29 00A75B29 00A65A29 00A65828
00A55728 00A45628 00A45528 00A35428
00A35328 00A25128 00A25028 00A14F28
00A04E27 00A04D27 009F4C27 009F4A27
009E4927 009E4827 009D4727 009C4627
009C4427 009B4326 009B4226 009A4126
009A4026 00993F26 00993D26 00983C26
00973B26 00973A26 00963925 00963825
00953625 00953525 00943425 00E2EBFE
00E1EAFE 00E1E9FE 00E0E8FE 00DFE7FE
00DEE6FE 00DEE5FE 00DDE4FE 00DCE3FE
00DBE2FE 00DBE1FD 00DAE0FD 00D9DFFD
00D8DEFD 00D8DDFD 00D7DCFD 00D6DBFD
00D6DAFD 00D5D9FD 00D4D8FD 00D3D7FD
00D3D6FD 00D2D5FD 00D1D4FD 00D0D3FD
00D0D2FD 00CFD1FD 00CED0FD 00CED0FD
00CDCEFC 00CCCDFC 00CBCCFC 00CACBFC
00CACBFC 00C9C9FC 00C8C8FC 00C8C7FC
00C7C6FC 00C6C5FC 00C5C4FC 00C4C3FC
00C4C2FC 00C3C1FC 00C2C0FC 00C1BFFC
00C1BEFC 00C0BDFC 00BFBCFB 00BEBBFB
00BEBAFB 00BDB9FB 00BCB8FB 00BBB7FB
00BBB6FB 00BAB5FB 00B9B4FB 00B9B3FB
00B8B2FB 00B8B1FB 00B8B0FB 00B7AFFB
00B7AEFB 00B7ADFB 00B6ABFB 00B6AAFA
00B6A9FA 00B5A8FA 00B5A7FA 00B5A6FA
00B4A5FA 00B4A4FA 00B3A3FA 00B3A1FA
00B3A0FA 00B29FFA 00B29EFA 00B29DFA
00B19CFA 00B19BFA 00B19AFA 00B098FA
00B097F9 00B096F9 00AF95F9 00AF94F9
00AE93F9 00AE91F9 00AE90F9 00AD8FF9
00AD8EF9 00AD8DF9 00AC8BF9 00AC8AF9
00AB89F9 00AB88F9 00AB87F9 00AA85F9
00AA84F8 00AA83F8 00A982F8 00A980F8
00A87FF8 00A87EF8 00A87DF8 00A77BF8
00A77AF8 00A679F8 00A678F8 00A676F8
00A575F8 00A574F8 00A472F8 00A471F7
00A370F7 00A36EF7 00A36DF7 00A26BF7
00A26AF7 00A169F7 00A167F7 00A166F6
00A066F5 00A065F5 00A064F4 009F63F4
009F62F3 009F61F2 009F60F2 009E5FF1
009E5EF0 009E5DF0 009D5CEF 009D5BEE
009D5AEE 009C59ED 009C58ED 009C57EC
009C56EB 009B55EB 009B54EA 009B53E9
009A52E9 009A51E8 009A50E7 009A4FE7
00994EE6 00994DE5 00994CE5 00984BE4
00984AE3 009849E3 009748E2 009747E1
009746E1 009645E0 009644DF 009642DF
009541DE 009540DD 00953FDD 00953EDC
00943DDB 00943CDA 00943BDA 00933AD9
009339D8 009338D8 009237D7 009235D6
009234D5 009133D5 009132D4 009131D3
009030D3 00902FD2 00902ED1 008F2CD0
008F2BD0 008E2ACF 008E29CE 008E28CD
008D26CC 008D25CC 008D24CB 008C23CA
008C22C9 008C20C8 008B1FC8 008B1EC7
008A1CC6 008A1BC5 008A1BC4 00891AC3
00891AC2 008919C1 008919BF 008819BE
008818BD 008818BC 008717BB 008717BA
008717B8 008616B7 008616B6 008615B5
008615B4 008515B3 008514B1 008514B0
008413AF 008413AE 008413AD 008412AC
008312AA 008311A9 008311A8 008211A7
008210A6 008210A5 00810FA3 00810FA2
00810FA1 00810EA0 00800E9F 00800D9E
00800D9C 007F0D9B 007F0C9A 007F0C99
007F0B98 007E0B97 007E0B95 007E0A94
007D0A93 007D0992 007D0991 007C0990
007C088F 007C088D 007C078C 007B078B
007B078A 007B0689 007A0688 007A0586
007A0585 007A0584 00790483 00790482
00790381 00780380 0078037E 0078027D
0078027C 0077017B 0077017A 0087080D
00880811 00890815 008A0818 008A081B
008B081E 008C0821 008C0824 008D0826
008E0829 008E082B 008F082E 008F0830
00900832 00900835 00910837 00910839
0092083B 0092083D 0093083F 00930841
00940843 00940845 00950847 00950849
0096084B 0096094D 0097094F 00970951
00980953 00980954 00980956 00990958
0099095A 009A095C 009A095D 009B095F
009B0961 009B0963 009C0964 009C0966
009D0968 009D0969 009D096B 009E096D
009E096F 009F0970 009F0972 009F0974
00A00975 00A00977 00A10979 00A1097A
00A1097C 00A2097E 00A2097F 00A30981
00A30982 00A30984 00A40986 00A40987
00A50989 00A5098B 00A40A8C 00A30C8E
00A10E90 00A01092 009F1293 009D1395
009C1597 009B1798 009A189A 00991A9B
00981B9C 00971D9E 00961E9F 00951FA1
009321A2 009222A3 009223A5 009125A6
009026A7 008F27A8 008E29AA 008D2AAB
008C2BAC 008B2CAD 008A2EAE 00892FAF
008830B1 008731B2 008732B3 008634B4
008535B5 008436B6 008337B7 008238B8
008139BA 00813ABB 00803CBC 007F3DBD
007E3EBE 007D3FBF 007D40C0 007C41C1
007B42C2 007A43C3 007944C4 007945C5
007846C6 007747C7 007649C8 00764AC9
00754BCA 00744CCB 00734DCC 00724ECD
00724FCE 007150CF 007051D0 006F52D1
006F53D2 006E54D3 006D55D4 006D56D5
006C57D6 006B58D7 006A59D8 006A5AD9
00695BDA 00685CDB 00675DDB 00665FDC
006560DD 006561DD 006463DE 006364DE
006265DF 006167DF 006068E0 006069E0
005F6BE1 005E6CE1 005D6DE2 005C6FE2
005C70E2 005B71E3 005A73E3 005974E4
005875E4 005876E5 005778E5 005679E6
00557AE6 00547BE7 00547DE7 00537EE8
00527FE8 005180E9 005181E9 005083E9
004F84EA 004E85EA 004E86EB 004D88EB
004C89EC 004B8AEC 004B8BED 004A8CED
00498DEE 00488FEE 004890EE 004791EF
004692EF 004593F0 004595F0 004496F1
004397F1 004298F2 004299F2 00419AF2
00409CF3 00409DF3 003F9EF4 003E9FF4
003DA0F5 003DA1F5 003CA2F5 003BA4F6
003BA5F6 003AA6F7 0039A7F7 0038A8F8
0038A9F8 0037AAF8 0036ACF9 0036ADF9
0035AEFA 0034AFFA 0033B0FB 0033B1FB
0032B2FB 0031B4FC 0031B5FC 0030B6FD
002FB7FD 002EB8FE 002EB9FE 002DBAFE
002CBBFF 002CBDFF 002CBEFE 002BC0FE
002BC1FE 002BC2FD 002BC4FD 002AC5FD
002AC7FC 002AC8FC 002AC9FC 0029CBFB
0029CCFB 0029CEFB 0029CFFA 0028D0FA
0028D2FA 0028D3F9 0028D4F9 0027D6F9
0027D7F8 0027D8F8 0027DAF8 0026DBF7
0026DDF7 0026DEF7 0026DFF6 0025E0F6
0025E2F6 0025E3F5 0025E4F5 0024E6F5
0024E7F4 0024E8F4 0024EAF4 0024EBF3
0023ECF3 0023EEF3 0023EFF3 0023F0F2
0022F1F2 0022F3F2 0022F4F1 0022F5F1
0021F6F1 0021F8F0 0021F9F0 000000FF
000006FF 00000CFF 000012FF 000018FF
00001EFF 000024FF 00002AFF 000030FF
000036FF 00003CFF 000042FF 000048FF
00004EFF 000054FF 00005AFF 000060FF
000066FF 00006CFF 000072FF 000078FF
00007EFF 000084FF 00008AFF 000090FF
000096FF 00009CFF 0000A2FF 0000A8FF
0000AEFF 0000B4FF 0000BAFF 0000C0FF
0000C6FF 0000CCFF 0000D2FF 0000D8FF
0000DEFF 0000E4FF 0000EAFF 0000F0FF
0000F6FF 0000FCFF 0000FFFC 0000FFF6
0000FFF0 0000FFEA 0000FFE4 0000FFDE
0000FFD8 0000FFD2 0000FFCC 0000FFC6
0000FFC0 0000FFBA 0000FFB4 0000FFAE
0000FFA8 0000FFA2 0000FF9C 0000FF96
0000FF90 0000FF8A 0000FF84 0000FF7E
0000FF78 0000FF72 0000FF6C 0000FF66
0000FF60 0000FF5A 0000FF54 0000FF4E
0000FF48 0000FF42 0000FF3C 0000FF36
0000FF30 0000FF2A 0000FF24 0000FF1E
0000FF18 0000FF12 0000FF0C 0000FF06
0000FF00 0006FF00 000CFF00 0012FF00
0018FF00 001EFF00 0024FF00 002AFF00
0030FF00 0036FF00 003CFF00 0042FF00
0048FF00 004EFF00 0054FF00 005AFF00
0060FF00 0066FF00 006CFF00 0072FF00
0078FF00 007EFF00 0084FF00 008AFF00
0090FF00 0096FF00 009CFF00 00A2FF00
00A8FF00 00AEFF00 00B4FF00 00BAFF00
00C0FF00 00C6FF00 00CCFF00 00D2FF00
00D8FF00 00DEFF00 00E4FF00 00EAFF00
00F0FF00 00F6FF00 00FCFF00 00FFFC00
00FFF600 00FFF000 00FFEA00 00FFE400
00FFDE00 00FFD800 00FFD200 00FFCC00
00FFC600 00FFC000 00FFBA00 00FFB400
00FFAE00 00FFA800 00FFA200 00FF9C00
00FF9600 00FF9000 00FF8A00 00FF8400
00FF7E00 00FF7800 00FF7200 00FF6C00
00FF6600 00FF6000 00FF5A00 00FF5400
00FF4E00 00FF4800 00FF4200 00FF3C00
00FF3600 00FF3000 00FF2A00 00FF2400
00FF1E00 00FF1800 00FF1200 00FF0C00
00FF0600 00FF0000 00FF0006 00FF000C
00FF0012 00FF0018 00FF001E 00FF0024
00FF002A 00FF0030 00FF0036 00FF003C
00FF0042 00FF0048 00FF004E 00FF0054
00FF005A 00FF0060 00FF0066 00FF006C
00FF0072 00FF0078 00FF007E 00FF0084
00FF008A 00FF0090 00FF0096 00FF009C
00FF00A2 00FF00A8 00FF00AE 00FF00B4
00FF00BA 00FF00C0 00FF00C6 00FF00CC
00FF00D2 00FF00D8 00FF00DE 00FF00E4
00FF00EA 00FF00F0 00FF00F6 00FF00FC
00FC00FF 00F600FF 00F000FF 00EA00FF
00E400FF 00DE00FF 00D800FF 00D200FF
00CC00FF 00C600FF 00C000FF 00BA00FF
00B400FF 00AE00FF 00A800FF 00A200FF
009C00FF 009600FF 009000FF 008A00FF
008400FF 007F00FE 007900FE 007300FE
006D00FE 006700FE 006100FE 005B00FE
005500FE 004F00FE 004900FE 004300FE
003D00FE 003700FE 003100FE 002B00FE
002500FE 001F00FE 001900FE 001300FE
000D00FE 000700FE 000100FE
@00000B17
00000014 00000000 00527A03 01017C01
07020D1B 00000001 00000010 0000001C
FFFFD384 00000018 00000000
@00000B22
80010004 80000000 FCA3999A FA03999A
